/*

Copyright (c) 2015-2020 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * si5341_i2c_init
 */
module si5341_i2c_init (
    input  wire        clk,
    input  wire        rst,

    /*
     * I2C master interface
     */
    output wire [6:0]  cmd_address,
    output wire        cmd_start,
    output wire        cmd_read,
    output wire        cmd_write,
    output wire        cmd_write_multiple,
    output wire        cmd_stop,
    output wire        cmd_valid,
    input  wire        cmd_ready,

    output wire [7:0]  data_out,
    output wire        data_out_valid,
    input  wire        data_out_ready,
    output wire        data_out_last,

    /*
     * Status
     */
    output wire        busy,

    /*
     * Configuration
     */
    input  wire        start
);

/*

Generic module for I2C bus initialization.  Good for use when multiple devices
on an I2C bus must be initialized on system start without intervention of a
general-purpose processor.

Copy this file and change init_data and INIT_DATA_LEN as needed.

This module can be used in two modes: simple device initalization, or multiple
device initialization.  In multiple device mode, the same initialization sequence
can be performed on multiple different device addresses.  

To use single device mode, only use the start write to address and write data commands.
The module will generate the I2C commands in sequential order.  Terminate the list
with a 0 entry.  

To use the multiple device mode, use the start data and start address block commands
to set up lists of initialization data and device addresses.  The module enters
multiple device mode upon seeing a start data block command.  The module stores the
offset of the start of the data block and then skips ahead until it reaches a start
address block command.  The module will store the offset to the address block and
read the first address in the block.  Then it will jump back to the data block
and execute it, substituting the stored address for each current address write
command.  Upon reaching the start address block command, the module will read out the
next address and start again at the top of the data block.  If the module encounters
a start data block command while looking for an address, then it will store a new data
offset and then look for a start address block command.  Terminate the list with a 0
entry.  Normal address commands will operate normally inside a data block.

Commands:

00 0000000 : stop
00 0000001 : exit multiple device mode
00 0000011 : start write to current address
00 0001000 : start address block
00 0001001 : start data block
00 1000001 : send I2C stop
01 aaaaaaa : start write to address
1 dddddddd : write 8-bit data

Examples

write 0x11223344 to register 0x0004 on device at 0x50

01 1010000  start write to 0x50
1 00000000  write address 0x0004
1 00000100
1 00010001  write data 0x11223344
1 00100010
1 00110011
1 01000100
0 00000000  stop

write 0x11223344 to register 0x0004 on devices at 0x50, 0x51, 0x52, and 0x53

00 0001001  start data block
00 0000011  start write to current address
1 00000100
1 00010001  write data 0x11223344
1 00100010
1 00110011
1 01000100
00 0001000  start address block
01 1010000  address 0x50
01 1010000  address 0x51
01 1010000  address 0x52
01 1010000  address 0x53
00 0000000  stop

*/

// init_data ROM
localparam INIT_DATA_LEN = 2329;

reg [8:0] init_data [INIT_DATA_LEN-1:0];

initial begin
    // Select Mux
    init_data[0] = {2'b01, 7'h74};
    init_data[1] = {1'b1,  8'h00};
    init_data[2] = 9'd0;                // Stop
    init_data[3] = {2'b01, 7'h75};
    init_data[4] = {1'b1,  8'h02};
    init_data[5] = 9'd0;                // Stop

    init_data[6] = 9'b111111111;        // Delay 300ms

    // Commands From ClockBuildPro
    init_data[7] = {2'b01, 7'h77};
    init_data[8] = {1'b1,  8'h01};
    init_data[9] = {1'b1,  8'h0B};
    init_data[10] = {2'b01, 7'h77};
    init_data[11] = {1'b1,  8'h24};
    init_data[12] = {1'b1,  8'hC0};
    init_data[13] = {2'b01, 7'h77};
    init_data[14] = {1'b1,  8'h01};
    init_data[15] = {1'b1,  8'h0B};
    init_data[16] = {2'b01, 7'h77};
    init_data[17] = {1'b1,  8'h25};
    init_data[18] = {1'b1,  8'h00};
    init_data[19] = {2'b01, 7'h77};
    init_data[20] = {1'b1,  8'h01};
    init_data[21] = {1'b1,  8'h05};
    init_data[22] = {2'b01, 7'h77};
    init_data[23] = {1'b1,  8'h02};
    init_data[24] = {1'b1,  8'h01};
    init_data[25] = {2'b01, 7'h77};
    init_data[26] = {1'b1,  8'h01};
    init_data[27] = {1'b1,  8'h05};
    init_data[28] = {2'b01, 7'h77};
    init_data[29] = {1'b1,  8'h05};
    init_data[30] = {1'b1,  8'h03};
    init_data[31] = {2'b01, 7'h77};
    init_data[32] = {1'b1,  8'h01};
    init_data[33] = {1'b1,  8'h09};
    init_data[34] = {2'b01, 7'h77};
    init_data[35] = {1'b1,  8'h57};
    init_data[36] = {1'b1,  8'h17};
    init_data[37] = {2'b01, 7'h77};
    init_data[38] = {1'b1,  8'h01};
    init_data[39] = {1'b1,  8'h0B};
    init_data[40] = {2'b01, 7'h77};
    init_data[41] = {1'b1,  8'h4E};
    init_data[42] = {1'b1,  8'h1A};
 /*
    # End configuration preamble
    #
    # Delay 300 msec
    #    Delay is worst case time for device to complete any calibration
    #    that is running due to device state change previous to this script
    #    being processed.
    #
    # Start configuration registers
  */
    init_data[43] = {2'b01, 7'h77};
    init_data[44] = {1'b1,  8'h01};
    init_data[45] = {1'b1,  8'h00};
    init_data[46] = {2'b01, 7'h77};
    init_data[47] = {1'b1,  8'h06};
    init_data[48] = {1'b1,  8'h00};
    init_data[49] = {2'b01, 7'h77};
    init_data[50] = {1'b1,  8'h01};
    init_data[51] = {1'b1,  8'h00};
    init_data[52] = {2'b01, 7'h77};
    init_data[53] = {1'b1,  8'h07};
    init_data[54] = {1'b1,  8'h00};
    init_data[55] = {2'b01, 7'h77};
    init_data[56] = {1'b1,  8'h01};
    init_data[57] = {1'b1,  8'h00};
    init_data[58] = {2'b01, 7'h77};
    init_data[59] = {1'b1,  8'h08};
    init_data[60] = {1'b1,  8'h00};
    init_data[61] = {2'b01, 7'h77};
    init_data[62] = {1'b1,  8'h01};
    init_data[63] = {1'b1,  8'h00};
    init_data[64] = {2'b01, 7'h77};
    init_data[65] = {1'b1,  8'h0B};
    init_data[66] = {1'b1,  8'h74};
    init_data[67] = {2'b01, 7'h77};
    init_data[68] = {1'b1,  8'h01};
    init_data[69] = {1'b1,  8'h00};
    init_data[70] = {2'b01, 7'h77};
    init_data[71] = {1'b1,  8'h17};
    init_data[72] = {1'b1,  8'hD0};
    init_data[73] = {2'b01, 7'h77};
    init_data[74] = {1'b1,  8'h01};
    init_data[75] = {1'b1,  8'h00};
    init_data[76] = {2'b01, 7'h77};
    init_data[77] = {1'b1,  8'h18};
    init_data[78] = {1'b1,  8'hFE};
    init_data[79] = {2'b01, 7'h77};
    init_data[80] = {1'b1,  8'h01};
    init_data[81] = {1'b1,  8'h00};
    init_data[82] = {2'b01, 7'h77};
    init_data[83] = {1'b1,  8'h21};
    init_data[84] = {1'b1,  8'h09};
    init_data[85] = {2'b01, 7'h77};
    init_data[86] = {1'b1,  8'h01};
    init_data[87] = {1'b1,  8'h00};
    init_data[88] = {2'b01, 7'h77};
    init_data[89] = {1'b1,  8'h22};
    init_data[90] = {1'b1,  8'h00};
    init_data[91] = {2'b01, 7'h77};
    init_data[92] = {1'b1,  8'h01};
    init_data[93] = {1'b1,  8'h00};
    init_data[94] = {2'b01, 7'h77};
    init_data[95] = {1'b1,  8'h2B};
    init_data[96] = {1'b1,  8'h02};
    init_data[97] = {2'b01, 7'h77};
    init_data[98] = {1'b1,  8'h01};
    init_data[99] = {1'b1,  8'h00};
    init_data[100] = {2'b01, 7'h77};
    init_data[101] = {1'b1,  8'h2C};
    init_data[102] = {1'b1,  8'h31};
    init_data[103] = {2'b01, 7'h77};
    init_data[104] = {1'b1,  8'h01};
    init_data[105] = {1'b1,  8'h00};
    init_data[106] = {2'b01, 7'h77};
    init_data[107] = {1'b1,  8'h2D};
    init_data[108] = {1'b1,  8'h01};
    init_data[109] = {2'b01, 7'h77};
    init_data[110] = {1'b1,  8'h01};
    init_data[111] = {1'b1,  8'h00};
    init_data[112] = {2'b01, 7'h77};
    init_data[113] = {1'b1,  8'h2E};
    init_data[114] = {1'b1,  8'hAE};
    init_data[115] = {2'b01, 7'h77};
    init_data[116] = {1'b1,  8'h01};
    init_data[117] = {1'b1,  8'h00};
    init_data[118] = {2'b01, 7'h77};
    init_data[119] = {1'b1,  8'h2F};
    init_data[120] = {1'b1,  8'h00};
    init_data[121] = {2'b01, 7'h77};
    init_data[122] = {1'b1,  8'h01};
    init_data[123] = {1'b1,  8'h00};
    init_data[124] = {2'b01, 7'h77};
    init_data[125] = {1'b1,  8'h30};
    init_data[126] = {1'b1,  8'h00};
    init_data[127] = {2'b01, 7'h77};
    init_data[128] = {1'b1,  8'h01};
    init_data[129] = {1'b1,  8'h00};
    init_data[130] = {2'b01, 7'h77};
    init_data[131] = {1'b1,  8'h31};
    init_data[132] = {1'b1,  8'h00};
    init_data[133] = {2'b01, 7'h77};
    init_data[134] = {1'b1,  8'h01};
    init_data[135] = {1'b1,  8'h00};
    init_data[136] = {2'b01, 7'h77};
    init_data[137] = {1'b1,  8'h32};
    init_data[138] = {1'b1,  8'h00};
    init_data[139] = {2'b01, 7'h77};
    init_data[140] = {1'b1,  8'h01};
    init_data[141] = {1'b1,  8'h00};
    init_data[142] = {2'b01, 7'h77};
    init_data[143] = {1'b1,  8'h33};
    init_data[144] = {1'b1,  8'h00};
    init_data[145] = {2'b01, 7'h77};
    init_data[146] = {1'b1,  8'h01};
    init_data[147] = {1'b1,  8'h00};
    init_data[148] = {2'b01, 7'h77};
    init_data[149] = {1'b1,  8'h34};
    init_data[150] = {1'b1,  8'h00};
    init_data[151] = {2'b01, 7'h77};
    init_data[152] = {1'b1,  8'h01};
    init_data[153] = {1'b1,  8'h00};
    init_data[154] = {2'b01, 7'h77};
    init_data[155] = {1'b1,  8'h35};
    init_data[156] = {1'b1,  8'h00};
    init_data[157] = {2'b01, 7'h77};
    init_data[158] = {1'b1,  8'h01};
    init_data[159] = {1'b1,  8'h00};
    init_data[160] = {2'b01, 7'h77};
    init_data[161] = {1'b1,  8'h36};
    init_data[162] = {1'b1,  8'hAE};
    init_data[163] = {2'b01, 7'h77};
    init_data[164] = {1'b1,  8'h01};
    init_data[165] = {1'b1,  8'h00};
    init_data[166] = {2'b01, 7'h77};
    init_data[167] = {1'b1,  8'h37};
    init_data[168] = {1'b1,  8'h00};
    init_data[169] = {2'b01, 7'h77};
    init_data[170] = {1'b1,  8'h01};
    init_data[171] = {1'b1,  8'h00};
    init_data[172] = {2'b01, 7'h77};
    init_data[173] = {1'b1,  8'h38};
    init_data[174] = {1'b1,  8'h00};
    init_data[175] = {2'b01, 7'h77};
    init_data[176] = {1'b1,  8'h01};
    init_data[177] = {1'b1,  8'h00};
    init_data[178] = {2'b01, 7'h77};
    init_data[179] = {1'b1,  8'h39};
    init_data[180] = {1'b1,  8'h00};
    init_data[181] = {2'b01, 7'h77};
    init_data[182] = {1'b1,  8'h01};
    init_data[183] = {1'b1,  8'h00};
    init_data[184] = {2'b01, 7'h77};
    init_data[185] = {1'b1,  8'h3A};
    init_data[186] = {1'b1,  8'h00};
    init_data[187] = {2'b01, 7'h77};
    init_data[188] = {1'b1,  8'h01};
    init_data[189] = {1'b1,  8'h00};
    init_data[190] = {2'b01, 7'h77};
    init_data[191] = {1'b1,  8'h3B};
    init_data[192] = {1'b1,  8'h00};
    init_data[193] = {2'b01, 7'h77};
    init_data[194] = {1'b1,  8'h01};
    init_data[195] = {1'b1,  8'h00};
    init_data[196] = {2'b01, 7'h77};
    init_data[197] = {1'b1,  8'h3C};
    init_data[198] = {1'b1,  8'h00};
    init_data[199] = {2'b01, 7'h77};
    init_data[200] = {1'b1,  8'h01};
    init_data[201] = {1'b1,  8'h00};
    init_data[202] = {2'b01, 7'h77};
    init_data[203] = {1'b1,  8'h3D};
    init_data[204] = {1'b1,  8'h00};
    init_data[205] = {2'b01, 7'h77};
    init_data[206] = {1'b1,  8'h01};
    init_data[207] = {1'b1,  8'h00};
    init_data[208] = {2'b01, 7'h77};
    init_data[209] = {1'b1,  8'h41};
    init_data[210] = {1'b1,  8'h07};
    init_data[211] = {2'b01, 7'h77};
    init_data[212] = {1'b1,  8'h01};
    init_data[213] = {1'b1,  8'h00};
    init_data[214] = {2'b01, 7'h77};
    init_data[215] = {1'b1,  8'h42};
    init_data[216] = {1'b1,  8'h00};
    init_data[217] = {2'b01, 7'h77};
    init_data[218] = {1'b1,  8'h01};
    init_data[219] = {1'b1,  8'h00};
    init_data[220] = {2'b01, 7'h77};
    init_data[221] = {1'b1,  8'h43};
    init_data[222] = {1'b1,  8'h00};
    init_data[223] = {2'b01, 7'h77};
    init_data[224] = {1'b1,  8'h01};
    init_data[225] = {1'b1,  8'h00};
    init_data[226] = {2'b01, 7'h77};
    init_data[227] = {1'b1,  8'h44};
    init_data[228] = {1'b1,  8'h00};
    init_data[229] = {2'b01, 7'h77};
    init_data[230] = {1'b1,  8'h01};
    init_data[231] = {1'b1,  8'h00};
    init_data[232] = {2'b01, 7'h77};
    init_data[233] = {1'b1,  8'h9E};
    init_data[234] = {1'b1,  8'h00};
    init_data[235] = {2'b01, 7'h77};
    init_data[236] = {1'b1,  8'h01};
    init_data[237] = {1'b1,  8'h01};
    init_data[238] = {2'b01, 7'h77};
    init_data[239] = {1'b1,  8'h02};
    init_data[240] = {1'b1,  8'h01};
    init_data[241] = {2'b01, 7'h77};
    init_data[242] = {1'b1,  8'h01};
    init_data[243] = {1'b1,  8'h01};
    init_data[244] = {2'b01, 7'h77};
    init_data[245] = {1'b1,  8'h08};
    init_data[246] = {1'b1,  8'h06};
    init_data[247] = {2'b01, 7'h77};
    init_data[248] = {1'b1,  8'h01};
    init_data[249] = {1'b1,  8'h01};
    init_data[250] = {2'b01, 7'h77};
    init_data[251] = {1'b1,  8'h09};
    init_data[252] = {1'b1,  8'h09};
    init_data[253] = {2'b01, 7'h77};
    init_data[254] = {1'b1,  8'h01};
    init_data[255] = {1'b1,  8'h01};
    init_data[256] = {2'b01, 7'h77};
    init_data[257] = {1'b1,  8'h0A};
    init_data[258] = {1'b1,  8'h33};
    init_data[259] = {2'b01, 7'h77};
    init_data[260] = {1'b1,  8'h01};
    init_data[261] = {1'b1,  8'h01};
    init_data[262] = {2'b01, 7'h77};
    init_data[263] = {1'b1,  8'h0B};
    init_data[264] = {1'b1,  8'h08};
    init_data[265] = {2'b01, 7'h77};
    init_data[266] = {1'b1,  8'h01};
    init_data[267] = {1'b1,  8'h01};
    init_data[268] = {2'b01, 7'h77};
    init_data[269] = {1'b1,  8'h0D};
    init_data[270] = {1'b1,  8'h06};
    init_data[271] = {2'b01, 7'h77};
    init_data[272] = {1'b1,  8'h01};
    init_data[273] = {1'b1,  8'h01};
    init_data[274] = {2'b01, 7'h77};
    init_data[275] = {1'b1,  8'h0E};
    init_data[276] = {1'b1,  8'h09};
    init_data[277] = {2'b01, 7'h77};
    init_data[278] = {1'b1,  8'h01};
    init_data[279] = {1'b1,  8'h01};
    init_data[280] = {2'b01, 7'h77};
    init_data[281] = {1'b1,  8'h0F};
    init_data[282] = {1'b1,  8'h33};
    init_data[283] = {2'b01, 7'h77};
    init_data[284] = {1'b1,  8'h01};
    init_data[285] = {1'b1,  8'h01};
    init_data[286] = {2'b01, 7'h77};
    init_data[287] = {1'b1,  8'h10};
    init_data[288] = {1'b1,  8'h08};
    init_data[289] = {2'b01, 7'h77};
    init_data[290] = {1'b1,  8'h01};
    init_data[291] = {1'b1,  8'h01};
    init_data[292] = {2'b01, 7'h77};
    init_data[293] = {1'b1,  8'h12};
    init_data[294] = {1'b1,  8'h06};
    init_data[295] = {2'b01, 7'h77};
    init_data[296] = {1'b1,  8'h01};
    init_data[297] = {1'b1,  8'h01};
    init_data[298] = {2'b01, 7'h77};
    init_data[299] = {1'b1,  8'h13};
    init_data[300] = {1'b1,  8'h09};
    init_data[301] = {2'b01, 7'h77};
    init_data[302] = {1'b1,  8'h01};
    init_data[303] = {1'b1,  8'h01};
    init_data[304] = {2'b01, 7'h77};
    init_data[305] = {1'b1,  8'h14};
    init_data[306] = {1'b1,  8'h33};
    init_data[307] = {2'b01, 7'h77};
    init_data[308] = {1'b1,  8'h01};
    init_data[309] = {1'b1,  8'h01};
    init_data[310] = {2'b01, 7'h77};
    init_data[311] = {1'b1,  8'h15};
    init_data[312] = {1'b1,  8'h08};
    init_data[313] = {2'b01, 7'h77};
    init_data[314] = {1'b1,  8'h01};
    init_data[315] = {1'b1,  8'h01};
    init_data[316] = {2'b01, 7'h77};
    init_data[317] = {1'b1,  8'h17};
    init_data[318] = {1'b1,  8'h06};
    init_data[319] = {2'b01, 7'h77};
    init_data[320] = {1'b1,  8'h01};
    init_data[321] = {1'b1,  8'h01};
    init_data[322] = {2'b01, 7'h77};
    init_data[323] = {1'b1,  8'h18};
    init_data[324] = {1'b1,  8'h09};
    init_data[325] = {2'b01, 7'h77};
    init_data[326] = {1'b1,  8'h01};
    init_data[327] = {1'b1,  8'h01};
    init_data[328] = {2'b01, 7'h77};
    init_data[329] = {1'b1,  8'h19};
    init_data[330] = {1'b1,  8'h33};
    init_data[331] = {2'b01, 7'h77};
    init_data[332] = {1'b1,  8'h01};
    init_data[333] = {1'b1,  8'h01};
    init_data[334] = {2'b01, 7'h77};
    init_data[335] = {1'b1,  8'h1A};
    init_data[336] = {1'b1,  8'h08};
    init_data[337] = {2'b01, 7'h77};
    init_data[338] = {1'b1,  8'h01};
    init_data[339] = {1'b1,  8'h01};
    init_data[340] = {2'b01, 7'h77};
    init_data[341] = {1'b1,  8'h1C};
    init_data[342] = {1'b1,  8'h06};
    init_data[343] = {2'b01, 7'h77};
    init_data[344] = {1'b1,  8'h01};
    init_data[345] = {1'b1,  8'h01};
    init_data[346] = {2'b01, 7'h77};
    init_data[347] = {1'b1,  8'h1D};
    init_data[348] = {1'b1,  8'h09};
    init_data[349] = {2'b01, 7'h77};
    init_data[350] = {1'b1,  8'h01};
    init_data[351] = {1'b1,  8'h01};
    init_data[352] = {2'b01, 7'h77};
    init_data[353] = {1'b1,  8'h1E};
    init_data[354] = {1'b1,  8'h33};
    init_data[355] = {2'b01, 7'h77};
    init_data[356] = {1'b1,  8'h01};
    init_data[357] = {1'b1,  8'h01};
    init_data[358] = {2'b01, 7'h77};
    init_data[359] = {1'b1,  8'h1F};
    init_data[360] = {1'b1,  8'h08};
    init_data[361] = {2'b01, 7'h77};
    init_data[362] = {1'b1,  8'h01};
    init_data[363] = {1'b1,  8'h01};
    init_data[364] = {2'b01, 7'h77};
    init_data[365] = {1'b1,  8'h21};
    init_data[366] = {1'b1,  8'h06};
    init_data[367] = {2'b01, 7'h77};
    init_data[368] = {1'b1,  8'h01};
    init_data[369] = {1'b1,  8'h01};
    init_data[370] = {2'b01, 7'h77};
    init_data[371] = {1'b1,  8'h22};
    init_data[372] = {1'b1,  8'h09};
    init_data[373] = {2'b01, 7'h77};
    init_data[374] = {1'b1,  8'h01};
    init_data[375] = {1'b1,  8'h01};
    init_data[376] = {2'b01, 7'h77};
    init_data[377] = {1'b1,  8'h23};
    init_data[378] = {1'b1,  8'h33};
    init_data[379] = {2'b01, 7'h77};
    init_data[380] = {1'b1,  8'h01};
    init_data[381] = {1'b1,  8'h01};
    init_data[382] = {2'b01, 7'h77};
    init_data[383] = {1'b1,  8'h24};
    init_data[384] = {1'b1,  8'h08};
    init_data[385] = {2'b01, 7'h77};
    init_data[386] = {1'b1,  8'h01};
    init_data[387] = {1'b1,  8'h01};
    init_data[388] = {2'b01, 7'h77};
    init_data[389] = {1'b1,  8'h26};
    init_data[390] = {1'b1,  8'h06};
    init_data[391] = {2'b01, 7'h77};
    init_data[392] = {1'b1,  8'h01};
    init_data[393] = {1'b1,  8'h01};
    init_data[394] = {2'b01, 7'h77};
    init_data[395] = {1'b1,  8'h27};
    init_data[396] = {1'b1,  8'h09};
    init_data[397] = {2'b01, 7'h77};
    init_data[398] = {1'b1,  8'h01};
    init_data[399] = {1'b1,  8'h01};
    init_data[400] = {2'b01, 7'h77};
    init_data[401] = {1'b1,  8'h28};
    init_data[402] = {1'b1,  8'h33};
    init_data[403] = {2'b01, 7'h77};
    init_data[404] = {1'b1,  8'h01};
    init_data[405] = {1'b1,  8'h01};
    init_data[406] = {2'b01, 7'h77};
    init_data[407] = {1'b1,  8'h29};
    init_data[408] = {1'b1,  8'h08};
    init_data[409] = {2'b01, 7'h77};
    init_data[410] = {1'b1,  8'h01};
    init_data[411] = {1'b1,  8'h01};
    init_data[412] = {2'b01, 7'h77};
    init_data[413] = {1'b1,  8'h2B};
    init_data[414] = {1'b1,  8'h06};
    init_data[415] = {2'b01, 7'h77};
    init_data[416] = {1'b1,  8'h01};
    init_data[417] = {1'b1,  8'h01};
    init_data[418] = {2'b01, 7'h77};
    init_data[419] = {1'b1,  8'h2C};
    init_data[420] = {1'b1,  8'h09};
    init_data[421] = {2'b01, 7'h77};
    init_data[422] = {1'b1,  8'h01};
    init_data[423] = {1'b1,  8'h01};
    init_data[424] = {2'b01, 7'h77};
    init_data[425] = {1'b1,  8'h2D};
    init_data[426] = {1'b1,  8'h33};
    init_data[427] = {2'b01, 7'h77};
    init_data[428] = {1'b1,  8'h01};
    init_data[429] = {1'b1,  8'h01};
    init_data[430] = {2'b01, 7'h77};
    init_data[431] = {1'b1,  8'h2E};
    init_data[432] = {1'b1,  8'h08};
    init_data[433] = {2'b01, 7'h77};
    init_data[434] = {1'b1,  8'h01};
    init_data[435] = {1'b1,  8'h01};
    init_data[436] = {2'b01, 7'h77};
    init_data[437] = {1'b1,  8'h30};
    init_data[438] = {1'b1,  8'h01};
    init_data[439] = {2'b01, 7'h77};
    init_data[440] = {1'b1,  8'h01};
    init_data[441] = {1'b1,  8'h01};
    init_data[442] = {2'b01, 7'h77};
    init_data[443] = {1'b1,  8'h31};
    init_data[444] = {1'b1,  8'h09};
    init_data[445] = {2'b01, 7'h77};
    init_data[446] = {1'b1,  8'h01};
    init_data[447] = {1'b1,  8'h01};
    init_data[448] = {2'b01, 7'h77};
    init_data[449] = {1'b1,  8'h32};
    init_data[450] = {1'b1,  8'h3B};
    init_data[451] = {2'b01, 7'h77};
    init_data[452] = {1'b1,  8'h01};
    init_data[453] = {1'b1,  8'h01};
    init_data[454] = {2'b01, 7'h77};
    init_data[455] = {1'b1,  8'h33};
    init_data[456] = {1'b1,  8'h28};
    init_data[457] = {2'b01, 7'h77};
    init_data[458] = {1'b1,  8'h01};
    init_data[459] = {1'b1,  8'h01};
    init_data[460] = {2'b01, 7'h77};
    init_data[461] = {1'b1,  8'h3A};
    init_data[462] = {1'b1,  8'h01};
    init_data[463] = {2'b01, 7'h77};
    init_data[464] = {1'b1,  8'h01};
    init_data[465] = {1'b1,  8'h01};
    init_data[466] = {2'b01, 7'h77};
    init_data[467] = {1'b1,  8'h3B};
    init_data[468] = {1'b1,  8'h09};
    init_data[469] = {2'b01, 7'h77};
    init_data[470] = {1'b1,  8'h01};
    init_data[471] = {1'b1,  8'h01};
    init_data[472] = {2'b01, 7'h77};
    init_data[473] = {1'b1,  8'h3C};
    init_data[474] = {1'b1,  8'h3B};
    init_data[475] = {2'b01, 7'h77};
    init_data[476] = {1'b1,  8'h01};
    init_data[477] = {1'b1,  8'h01};
    init_data[478] = {2'b01, 7'h77};
    init_data[479] = {1'b1,  8'h3D};
    init_data[480] = {1'b1,  8'h28};
    init_data[481] = {2'b01, 7'h77};
    init_data[482] = {1'b1,  8'h01};
    init_data[483] = {1'b1,  8'h01};
    init_data[484] = {2'b01, 7'h77};
    init_data[485] = {1'b1,  8'h3F};
    init_data[486] = {1'b1,  8'h00};
    init_data[487] = {2'b01, 7'h77};
    init_data[488] = {1'b1,  8'h01};
    init_data[489] = {1'b1,  8'h01};
    init_data[490] = {2'b01, 7'h77};
    init_data[491] = {1'b1,  8'h40};
    init_data[492] = {1'b1,  8'h00};
    init_data[493] = {2'b01, 7'h77};
    init_data[494] = {1'b1,  8'h01};
    init_data[495] = {1'b1,  8'h01};
    init_data[496] = {2'b01, 7'h77};
    init_data[497] = {1'b1,  8'h41};
    init_data[498] = {1'b1,  8'h40};
    init_data[499] = {2'b01, 7'h77};
    init_data[500] = {1'b1,  8'h01};
    init_data[501] = {1'b1,  8'h02};
    init_data[502] = {2'b01, 7'h77};
    init_data[503] = {1'b1,  8'h06};
    init_data[504] = {1'b1,  8'h00};
    init_data[505] = {2'b01, 7'h77};
    init_data[506] = {1'b1,  8'h01};
    init_data[507] = {1'b1,  8'h02};
    init_data[508] = {2'b01, 7'h77};
    init_data[509] = {1'b1,  8'h08};
    init_data[510] = {1'b1,  8'h02};
    init_data[511] = {2'b01, 7'h77};
    init_data[512] = {1'b1,  8'h01};
    init_data[513] = {1'b1,  8'h02};
    init_data[514] = {2'b01, 7'h77};
    init_data[515] = {1'b1,  8'h09};
    init_data[516] = {1'b1,  8'h00};
    init_data[517] = {2'b01, 7'h77};
    init_data[518] = {1'b1,  8'h01};
    init_data[519] = {1'b1,  8'h02};
    init_data[520] = {2'b01, 7'h77};
    init_data[521] = {1'b1,  8'h0A};
    init_data[522] = {1'b1,  8'h00};
    init_data[523] = {2'b01, 7'h77};
    init_data[524] = {1'b1,  8'h01};
    init_data[525] = {1'b1,  8'h02};
    init_data[526] = {2'b01, 7'h77};
    init_data[527] = {1'b1,  8'h0B};
    init_data[528] = {1'b1,  8'h00};
    init_data[529] = {2'b01, 7'h77};
    init_data[530] = {1'b1,  8'h01};
    init_data[531] = {1'b1,  8'h02};
    init_data[532] = {2'b01, 7'h77};
    init_data[533] = {1'b1,  8'h0C};
    init_data[534] = {1'b1,  8'h00};
    init_data[535] = {2'b01, 7'h77};
    init_data[536] = {1'b1,  8'h01};
    init_data[537] = {1'b1,  8'h02};
    init_data[538] = {2'b01, 7'h77};
    init_data[539] = {1'b1,  8'h0D};
    init_data[540] = {1'b1,  8'h00};
    init_data[541] = {2'b01, 7'h77};
    init_data[542] = {1'b1,  8'h01};
    init_data[543] = {1'b1,  8'h02};
    init_data[544] = {2'b01, 7'h77};
    init_data[545] = {1'b1,  8'h0E};
    init_data[546] = {1'b1,  8'h01};
    init_data[547] = {2'b01, 7'h77};
    init_data[548] = {1'b1,  8'h01};
    init_data[549] = {1'b1,  8'h02};
    init_data[550] = {2'b01, 7'h77};
    init_data[551] = {1'b1,  8'h0F};
    init_data[552] = {1'b1,  8'h00};
    init_data[553] = {2'b01, 7'h77};
    init_data[554] = {1'b1,  8'h01};
    init_data[555] = {1'b1,  8'h02};
    init_data[556] = {2'b01, 7'h77};
    init_data[557] = {1'b1,  8'h10};
    init_data[558] = {1'b1,  8'h00};
    init_data[559] = {2'b01, 7'h77};
    init_data[560] = {1'b1,  8'h01};
    init_data[561] = {1'b1,  8'h02};
    init_data[562] = {2'b01, 7'h77};
    init_data[563] = {1'b1,  8'h11};
    init_data[564] = {1'b1,  8'h00};
    init_data[565] = {2'b01, 7'h77};
    init_data[566] = {1'b1,  8'h01};
    init_data[567] = {1'b1,  8'h02};
    init_data[568] = {2'b01, 7'h77};
    init_data[569] = {1'b1,  8'h12};
    init_data[570] = {1'b1,  8'h00};
    init_data[571] = {2'b01, 7'h77};
    init_data[572] = {1'b1,  8'h01};
    init_data[573] = {1'b1,  8'h02};
    init_data[574] = {2'b01, 7'h77};
    init_data[575] = {1'b1,  8'h13};
    init_data[576] = {1'b1,  8'h00};
    init_data[577] = {2'b01, 7'h77};
    init_data[578] = {1'b1,  8'h01};
    init_data[579] = {1'b1,  8'h02};
    init_data[580] = {2'b01, 7'h77};
    init_data[581] = {1'b1,  8'h14};
    init_data[582] = {1'b1,  8'h00};
    init_data[583] = {2'b01, 7'h77};
    init_data[584] = {1'b1,  8'h01};
    init_data[585] = {1'b1,  8'h02};
    init_data[586] = {2'b01, 7'h77};
    init_data[587] = {1'b1,  8'h15};
    init_data[588] = {1'b1,  8'h00};
    init_data[589] = {2'b01, 7'h77};
    init_data[590] = {1'b1,  8'h01};
    init_data[591] = {1'b1,  8'h02};
    init_data[592] = {2'b01, 7'h77};
    init_data[593] = {1'b1,  8'h16};
    init_data[594] = {1'b1,  8'h00};
    init_data[595] = {2'b01, 7'h77};
    init_data[596] = {1'b1,  8'h01};
    init_data[597] = {1'b1,  8'h02};
    init_data[598] = {2'b01, 7'h77};
    init_data[599] = {1'b1,  8'h17};
    init_data[600] = {1'b1,  8'h00};
    init_data[601] = {2'b01, 7'h77};
    init_data[602] = {1'b1,  8'h01};
    init_data[603] = {1'b1,  8'h02};
    init_data[604] = {2'b01, 7'h77};
    init_data[605] = {1'b1,  8'h18};
    init_data[606] = {1'b1,  8'h00};
    init_data[607] = {2'b01, 7'h77};
    init_data[608] = {1'b1,  8'h01};
    init_data[609] = {1'b1,  8'h02};
    init_data[610] = {2'b01, 7'h77};
    init_data[611] = {1'b1,  8'h19};
    init_data[612] = {1'b1,  8'h00};
    init_data[613] = {2'b01, 7'h77};
    init_data[614] = {1'b1,  8'h01};
    init_data[615] = {1'b1,  8'h02};
    init_data[616] = {2'b01, 7'h77};
    init_data[617] = {1'b1,  8'h1A};
    init_data[618] = {1'b1,  8'h00};
    init_data[619] = {2'b01, 7'h77};
    init_data[620] = {1'b1,  8'h01};
    init_data[621] = {1'b1,  8'h02};
    init_data[622] = {2'b01, 7'h77};
    init_data[623] = {1'b1,  8'h1B};
    init_data[624] = {1'b1,  8'h00};
    init_data[625] = {2'b01, 7'h77};
    init_data[626] = {1'b1,  8'h01};
    init_data[627] = {1'b1,  8'h02};
    init_data[628] = {2'b01, 7'h77};
    init_data[629] = {1'b1,  8'h1C};
    init_data[630] = {1'b1,  8'h00};
    init_data[631] = {2'b01, 7'h77};
    init_data[632] = {1'b1,  8'h01};
    init_data[633] = {1'b1,  8'h02};
    init_data[634] = {2'b01, 7'h77};
    init_data[635] = {1'b1,  8'h1D};
    init_data[636] = {1'b1,  8'h00};
    init_data[637] = {2'b01, 7'h77};
    init_data[638] = {1'b1,  8'h01};
    init_data[639] = {1'b1,  8'h02};
    init_data[640] = {2'b01, 7'h77};
    init_data[641] = {1'b1,  8'h1E};
    init_data[642] = {1'b1,  8'h00};
    init_data[643] = {2'b01, 7'h77};
    init_data[644] = {1'b1,  8'h01};
    init_data[645] = {1'b1,  8'h02};
    init_data[646] = {2'b01, 7'h77};
    init_data[647] = {1'b1,  8'h1F};
    init_data[648] = {1'b1,  8'h00};
    init_data[649] = {2'b01, 7'h77};
    init_data[650] = {1'b1,  8'h01};
    init_data[651] = {1'b1,  8'h02};
    init_data[652] = {2'b01, 7'h77};
    init_data[653] = {1'b1,  8'h20};
    init_data[654] = {1'b1,  8'h00};
    init_data[655] = {2'b01, 7'h77};
    init_data[656] = {1'b1,  8'h01};
    init_data[657] = {1'b1,  8'h02};
    init_data[658] = {2'b01, 7'h77};
    init_data[659] = {1'b1,  8'h21};
    init_data[660] = {1'b1,  8'h00};
    init_data[661] = {2'b01, 7'h77};
    init_data[662] = {1'b1,  8'h01};
    init_data[663] = {1'b1,  8'h02};
    init_data[664] = {2'b01, 7'h77};
    init_data[665] = {1'b1,  8'h22};
    init_data[666] = {1'b1,  8'h00};
    init_data[667] = {2'b01, 7'h77};
    init_data[668] = {1'b1,  8'h01};
    init_data[669] = {1'b1,  8'h02};
    init_data[670] = {2'b01, 7'h77};
    init_data[671] = {1'b1,  8'h23};
    init_data[672] = {1'b1,  8'h00};
    init_data[673] = {2'b01, 7'h77};
    init_data[674] = {1'b1,  8'h01};
    init_data[675] = {1'b1,  8'h02};
    init_data[676] = {2'b01, 7'h77};
    init_data[677] = {1'b1,  8'h24};
    init_data[678] = {1'b1,  8'h00};
    init_data[679] = {2'b01, 7'h77};
    init_data[680] = {1'b1,  8'h01};
    init_data[681] = {1'b1,  8'h02};
    init_data[682] = {2'b01, 7'h77};
    init_data[683] = {1'b1,  8'h25};
    init_data[684] = {1'b1,  8'h00};
    init_data[685] = {2'b01, 7'h77};
    init_data[686] = {1'b1,  8'h01};
    init_data[687] = {1'b1,  8'h02};
    init_data[688] = {2'b01, 7'h77};
    init_data[689] = {1'b1,  8'h26};
    init_data[690] = {1'b1,  8'h00};
    init_data[691] = {2'b01, 7'h77};
    init_data[692] = {1'b1,  8'h01};
    init_data[693] = {1'b1,  8'h02};
    init_data[694] = {2'b01, 7'h77};
    init_data[695] = {1'b1,  8'h27};
    init_data[696] = {1'b1,  8'h00};
    init_data[697] = {2'b01, 7'h77};
    init_data[698] = {1'b1,  8'h01};
    init_data[699] = {1'b1,  8'h02};
    init_data[700] = {2'b01, 7'h77};
    init_data[701] = {1'b1,  8'h28};
    init_data[702] = {1'b1,  8'h00};
    init_data[703] = {2'b01, 7'h77};
    init_data[704] = {1'b1,  8'h01};
    init_data[705] = {1'b1,  8'h02};
    init_data[706] = {2'b01, 7'h77};
    init_data[707] = {1'b1,  8'h29};
    init_data[708] = {1'b1,  8'h00};
    init_data[709] = {2'b01, 7'h77};
    init_data[710] = {1'b1,  8'h01};
    init_data[711] = {1'b1,  8'h02};
    init_data[712] = {2'b01, 7'h77};
    init_data[713] = {1'b1,  8'h2A};
    init_data[714] = {1'b1,  8'h00};
    init_data[715] = {2'b01, 7'h77};
    init_data[716] = {1'b1,  8'h01};
    init_data[717] = {1'b1,  8'h02};
    init_data[718] = {2'b01, 7'h77};
    init_data[719] = {1'b1,  8'h2B};
    init_data[720] = {1'b1,  8'h00};
    init_data[721] = {2'b01, 7'h77};
    init_data[722] = {1'b1,  8'h01};
    init_data[723] = {1'b1,  8'h02};
    init_data[724] = {2'b01, 7'h77};
    init_data[725] = {1'b1,  8'h2C};
    init_data[726] = {1'b1,  8'h00};
    init_data[727] = {2'b01, 7'h77};
    init_data[728] = {1'b1,  8'h01};
    init_data[729] = {1'b1,  8'h02};
    init_data[730] = {2'b01, 7'h77};
    init_data[731] = {1'b1,  8'h2D};
    init_data[732] = {1'b1,  8'h00};
    init_data[733] = {2'b01, 7'h77};
    init_data[734] = {1'b1,  8'h01};
    init_data[735] = {1'b1,  8'h02};
    init_data[736] = {2'b01, 7'h77};
    init_data[737] = {1'b1,  8'h2E};
    init_data[738] = {1'b1,  8'h00};
    init_data[739] = {2'b01, 7'h77};
    init_data[740] = {1'b1,  8'h01};
    init_data[741] = {1'b1,  8'h02};
    init_data[742] = {2'b01, 7'h77};
    init_data[743] = {1'b1,  8'h2F};
    init_data[744] = {1'b1,  8'h00};
    init_data[745] = {2'b01, 7'h77};
    init_data[746] = {1'b1,  8'h01};
    init_data[747] = {1'b1,  8'h02};
    init_data[748] = {2'b01, 7'h77};
    init_data[749] = {1'b1,  8'h35};
    init_data[750] = {1'b1,  8'h00};
    init_data[751] = {2'b01, 7'h77};
    init_data[752] = {1'b1,  8'h01};
    init_data[753] = {1'b1,  8'h02};
    init_data[754] = {2'b01, 7'h77};
    init_data[755] = {1'b1,  8'h36};
    init_data[756] = {1'b1,  8'h00};
    init_data[757] = {2'b01, 7'h77};
    init_data[758] = {1'b1,  8'h01};
    init_data[759] = {1'b1,  8'h02};
    init_data[760] = {2'b01, 7'h77};
    init_data[761] = {1'b1,  8'h37};
    init_data[762] = {1'b1,  8'h00};
    init_data[763] = {2'b01, 7'h77};
    init_data[764] = {1'b1,  8'h01};
    init_data[765] = {1'b1,  8'h02};
    init_data[766] = {2'b01, 7'h77};
    init_data[767] = {1'b1,  8'h38};
    init_data[768] = {1'b1,  8'h90};
    init_data[769] = {2'b01, 7'h77};
    init_data[770] = {1'b1,  8'h01};
    init_data[771] = {1'b1,  8'h02};
    init_data[772] = {2'b01, 7'h77};
    init_data[773] = {1'b1,  8'h39};
    init_data[774] = {1'b1,  8'h54};
    init_data[775] = {2'b01, 7'h77};
    init_data[776] = {1'b1,  8'h01};
    init_data[777] = {1'b1,  8'h02};
    init_data[778] = {2'b01, 7'h77};
    init_data[779] = {1'b1,  8'h3A};
    init_data[780] = {1'b1,  8'h00};
    init_data[781] = {2'b01, 7'h77};
    init_data[782] = {1'b1,  8'h01};
    init_data[783] = {1'b1,  8'h02};
    init_data[784] = {2'b01, 7'h77};
    init_data[785] = {1'b1,  8'h3B};
    init_data[786] = {1'b1,  8'h00};
    init_data[787] = {2'b01, 7'h77};
    init_data[788] = {1'b1,  8'h01};
    init_data[789] = {1'b1,  8'h02};
    init_data[790] = {2'b01, 7'h77};
    init_data[791] = {1'b1,  8'h3C};
    init_data[792] = {1'b1,  8'h00};
    init_data[793] = {2'b01, 7'h77};
    init_data[794] = {1'b1,  8'h01};
    init_data[795] = {1'b1,  8'h02};
    init_data[796] = {2'b01, 7'h77};
    init_data[797] = {1'b1,  8'h3D};
    init_data[798] = {1'b1,  8'h00};
    init_data[799] = {2'b01, 7'h77};
    init_data[800] = {1'b1,  8'h01};
    init_data[801] = {1'b1,  8'h02};
    init_data[802] = {2'b01, 7'h77};
    init_data[803] = {1'b1,  8'h3E};
    init_data[804] = {1'b1,  8'h80};
    init_data[805] = {2'b01, 7'h77};
    init_data[806] = {1'b1,  8'h01};
    init_data[807] = {1'b1,  8'h02};
    init_data[808] = {2'b01, 7'h77};
    init_data[809] = {1'b1,  8'h4A};
    init_data[810] = {1'b1,  8'h00};
    init_data[811] = {2'b01, 7'h77};
    init_data[812] = {1'b1,  8'h01};
    init_data[813] = {1'b1,  8'h02};
    init_data[814] = {2'b01, 7'h77};
    init_data[815] = {1'b1,  8'h4B};
    init_data[816] = {1'b1,  8'h00};
    init_data[817] = {2'b01, 7'h77};
    init_data[818] = {1'b1,  8'h01};
    init_data[819] = {1'b1,  8'h02};
    init_data[820] = {2'b01, 7'h77};
    init_data[821] = {1'b1,  8'h4C};
    init_data[822] = {1'b1,  8'h00};
    init_data[823] = {2'b01, 7'h77};
    init_data[824] = {1'b1,  8'h01};
    init_data[825] = {1'b1,  8'h02};
    init_data[826] = {2'b01, 7'h77};
    init_data[827] = {1'b1,  8'h4D};
    init_data[828] = {1'b1,  8'h00};
    init_data[829] = {2'b01, 7'h77};
    init_data[830] = {1'b1,  8'h01};
    init_data[831] = {1'b1,  8'h02};
    init_data[832] = {2'b01, 7'h77};
    init_data[833] = {1'b1,  8'h4E};
    init_data[834] = {1'b1,  8'h00};
    init_data[835] = {2'b01, 7'h77};
    init_data[836] = {1'b1,  8'h01};
    init_data[837] = {1'b1,  8'h02};
    init_data[838] = {2'b01, 7'h77};
    init_data[839] = {1'b1,  8'h4F};
    init_data[840] = {1'b1,  8'h00};
    init_data[841] = {2'b01, 7'h77};
    init_data[842] = {1'b1,  8'h01};
    init_data[843] = {1'b1,  8'h02};
    init_data[844] = {2'b01, 7'h77};
    init_data[845] = {1'b1,  8'h50};
    init_data[846] = {1'b1,  8'h00};
    init_data[847] = {2'b01, 7'h77};
    init_data[848] = {1'b1,  8'h01};
    init_data[849] = {1'b1,  8'h02};
    init_data[850] = {2'b01, 7'h77};
    init_data[851] = {1'b1,  8'h51};
    init_data[852] = {1'b1,  8'h00};
    init_data[853] = {2'b01, 7'h77};
    init_data[854] = {1'b1,  8'h01};
    init_data[855] = {1'b1,  8'h02};
    init_data[856] = {2'b01, 7'h77};
    init_data[857] = {1'b1,  8'h52};
    init_data[858] = {1'b1,  8'h00};
    init_data[859] = {2'b01, 7'h77};
    init_data[860] = {1'b1,  8'h01};
    init_data[861] = {1'b1,  8'h02};
    init_data[862] = {2'b01, 7'h77};
    init_data[863] = {1'b1,  8'h53};
    init_data[864] = {1'b1,  8'h00};
    init_data[865] = {2'b01, 7'h77};
    init_data[866] = {1'b1,  8'h01};
    init_data[867] = {1'b1,  8'h02};
    init_data[868] = {2'b01, 7'h77};
    init_data[869] = {1'b1,  8'h54};
    init_data[870] = {1'b1,  8'h00};
    init_data[871] = {2'b01, 7'h77};
    init_data[872] = {1'b1,  8'h01};
    init_data[873] = {1'b1,  8'h02};
    init_data[874] = {2'b01, 7'h77};
    init_data[875] = {1'b1,  8'h55};
    init_data[876] = {1'b1,  8'h00};
    init_data[877] = {2'b01, 7'h77};
    init_data[878] = {1'b1,  8'h01};
    init_data[879] = {1'b1,  8'h02};
    init_data[880] = {2'b01, 7'h77};
    init_data[881] = {1'b1,  8'h56};
    init_data[882] = {1'b1,  8'h00};
    init_data[883] = {2'b01, 7'h77};
    init_data[884] = {1'b1,  8'h01};
    init_data[885] = {1'b1,  8'h02};
    init_data[886] = {2'b01, 7'h77};
    init_data[887] = {1'b1,  8'h57};
    init_data[888] = {1'b1,  8'h00};
    init_data[889] = {2'b01, 7'h77};
    init_data[890] = {1'b1,  8'h01};
    init_data[891] = {1'b1,  8'h02};
    init_data[892] = {2'b01, 7'h77};
    init_data[893] = {1'b1,  8'h58};
    init_data[894] = {1'b1,  8'h00};
    init_data[895] = {2'b01, 7'h77};
    init_data[896] = {1'b1,  8'h01};
    init_data[897] = {1'b1,  8'h02};
    init_data[898] = {2'b01, 7'h77};
    init_data[899] = {1'b1,  8'h59};
    init_data[900] = {1'b1,  8'h00};
    init_data[901] = {2'b01, 7'h77};
    init_data[902] = {1'b1,  8'h01};
    init_data[903] = {1'b1,  8'h02};
    init_data[904] = {2'b01, 7'h77};
    init_data[905] = {1'b1,  8'h5A};
    init_data[906] = {1'b1,  8'h00};
    init_data[907] = {2'b01, 7'h77};
    init_data[908] = {1'b1,  8'h01};
    init_data[909] = {1'b1,  8'h02};
    init_data[910] = {2'b01, 7'h77};
    init_data[911] = {1'b1,  8'h5B};
    init_data[912] = {1'b1,  8'h00};
    init_data[913] = {2'b01, 7'h77};
    init_data[914] = {1'b1,  8'h01};
    init_data[915] = {1'b1,  8'h02};
    init_data[916] = {2'b01, 7'h77};
    init_data[917] = {1'b1,  8'h5C};
    init_data[918] = {1'b1,  8'h00};
    init_data[919] = {2'b01, 7'h77};
    init_data[920] = {1'b1,  8'h01};
    init_data[921] = {1'b1,  8'h02};
    init_data[922] = {2'b01, 7'h77};
    init_data[923] = {1'b1,  8'h5D};
    init_data[924] = {1'b1,  8'h00};
    init_data[925] = {2'b01, 7'h77};
    init_data[926] = {1'b1,  8'h01};
    init_data[927] = {1'b1,  8'h02};
    init_data[928] = {2'b01, 7'h77};
    init_data[929] = {1'b1,  8'h5E};
    init_data[930] = {1'b1,  8'h00};
    init_data[931] = {2'b01, 7'h77};
    init_data[932] = {1'b1,  8'h01};
    init_data[933] = {1'b1,  8'h02};
    init_data[934] = {2'b01, 7'h77};
    init_data[935] = {1'b1,  8'h5F};
    init_data[936] = {1'b1,  8'h00};
    init_data[937] = {2'b01, 7'h77};
    init_data[938] = {1'b1,  8'h01};
    init_data[939] = {1'b1,  8'h02};
    init_data[940] = {2'b01, 7'h77};
    init_data[941] = {1'b1,  8'h60};
    init_data[942] = {1'b1,  8'h00};
    init_data[943] = {2'b01, 7'h77};
    init_data[944] = {1'b1,  8'h01};
    init_data[945] = {1'b1,  8'h02};
    init_data[946] = {2'b01, 7'h77};
    init_data[947] = {1'b1,  8'h61};
    init_data[948] = {1'b1,  8'h00};
    init_data[949] = {2'b01, 7'h77};
    init_data[950] = {1'b1,  8'h01};
    init_data[951] = {1'b1,  8'h02};
    init_data[952] = {2'b01, 7'h77};
    init_data[953] = {1'b1,  8'h62};
    init_data[954] = {1'b1,  8'h00};
    init_data[955] = {2'b01, 7'h77};
    init_data[956] = {1'b1,  8'h01};
    init_data[957] = {1'b1,  8'h02};
    init_data[958] = {2'b01, 7'h77};
    init_data[959] = {1'b1,  8'h63};
    init_data[960] = {1'b1,  8'h00};
    init_data[961] = {2'b01, 7'h77};
    init_data[962] = {1'b1,  8'h01};
    init_data[963] = {1'b1,  8'h02};
    init_data[964] = {2'b01, 7'h77};
    init_data[965] = {1'b1,  8'h64};
    init_data[966] = {1'b1,  8'h00};
    init_data[967] = {2'b01, 7'h77};
    init_data[968] = {1'b1,  8'h01};
    init_data[969] = {1'b1,  8'h02};
    init_data[970] = {2'b01, 7'h77};
    init_data[971] = {1'b1,  8'h68};
    init_data[972] = {1'b1,  8'h00};
    init_data[973] = {2'b01, 7'h77};
    init_data[974] = {1'b1,  8'h01};
    init_data[975] = {1'b1,  8'h02};
    init_data[976] = {2'b01, 7'h77};
    init_data[977] = {1'b1,  8'h69};
    init_data[978] = {1'b1,  8'h00};
    init_data[979] = {2'b01, 7'h77};
    init_data[980] = {1'b1,  8'h01};
    init_data[981] = {1'b1,  8'h02};
    init_data[982] = {2'b01, 7'h77};
    init_data[983] = {1'b1,  8'h6A};
    init_data[984] = {1'b1,  8'h00};
    init_data[985] = {2'b01, 7'h77};
    init_data[986] = {1'b1,  8'h01};
    init_data[987] = {1'b1,  8'h02};
    init_data[988] = {2'b01, 7'h77};
    init_data[989] = {1'b1,  8'h6B};
    init_data[990] = {1'b1,  8'h48};
    init_data[991] = {2'b01, 7'h77};
    init_data[992] = {1'b1,  8'h01};
    init_data[993] = {1'b1,  8'h02};
    init_data[994] = {2'b01, 7'h77};
    init_data[995] = {1'b1,  8'h6C};
    init_data[996] = {1'b1,  8'h54};
    init_data[997] = {2'b01, 7'h77};
    init_data[998] = {1'b1,  8'h01};
    init_data[999] = {1'b1,  8'h02};
    init_data[1000] = {2'b01, 7'h77};
    init_data[1001] = {1'b1,  8'h6D};
    init_data[1002] = {1'b1,  8'h47};
    init_data[1003] = {2'b01, 7'h77};
    init_data[1004] = {1'b1,  8'h01};
    init_data[1005] = {1'b1,  8'h02};
    init_data[1006] = {2'b01, 7'h77};
    init_data[1007] = {1'b1,  8'h6E};
    init_data[1008] = {1'b1,  8'h51};
    init_data[1009] = {2'b01, 7'h77};
    init_data[1010] = {1'b1,  8'h01};
    init_data[1011] = {1'b1,  8'h02};
    init_data[1012] = {2'b01, 7'h77};
    init_data[1013] = {1'b1,  8'h6F};
    init_data[1014] = {1'b1,  8'h53};
    init_data[1015] = {2'b01, 7'h77};
    init_data[1016] = {1'b1,  8'h01};
    init_data[1017] = {1'b1,  8'h02};
    init_data[1018] = {2'b01, 7'h77};
    init_data[1019] = {1'b1,  8'h70};
    init_data[1020] = {1'b1,  8'h46};
    init_data[1021] = {2'b01, 7'h77};
    init_data[1022] = {1'b1,  8'h01};
    init_data[1023] = {1'b1,  8'h02};
    init_data[1024] = {2'b01, 7'h77};
    init_data[1025] = {1'b1,  8'h71};
    init_data[1026] = {1'b1,  8'h50};
    init_data[1027] = {2'b01, 7'h77};
    init_data[1028] = {1'b1,  8'h01};
    init_data[1029] = {1'b1,  8'h02};
    init_data[1030] = {2'b01, 7'h77};
    init_data[1031] = {1'b1,  8'h72};
    init_data[1032] = {1'b1,  8'h00};
    init_data[1033] = {2'b01, 7'h77};
    init_data[1034] = {1'b1,  8'h01};
    init_data[1035] = {1'b1,  8'h03};
    init_data[1036] = {2'b01, 7'h77};
    init_data[1037] = {1'b1,  8'h02};
    init_data[1038] = {1'b1,  8'h00};
    init_data[1039] = {2'b01, 7'h77};
    init_data[1040] = {1'b1,  8'h01};
    init_data[1041] = {1'b1,  8'h03};
    init_data[1042] = {2'b01, 7'h77};
    init_data[1043] = {1'b1,  8'h03};
    init_data[1044] = {1'b1,  8'h00};
    init_data[1045] = {2'b01, 7'h77};
    init_data[1046] = {1'b1,  8'h01};
    init_data[1047] = {1'b1,  8'h03};
    init_data[1048] = {2'b01, 7'h77};
    init_data[1049] = {1'b1,  8'h04};
    init_data[1050] = {1'b1,  8'h00};
    init_data[1051] = {2'b01, 7'h77};
    init_data[1052] = {1'b1,  8'h01};
    init_data[1053] = {1'b1,  8'h03};
    init_data[1054] = {2'b01, 7'h77};
    init_data[1055] = {1'b1,  8'h05};
    init_data[1056] = {1'b1,  8'h80};
    init_data[1057] = {2'b01, 7'h77};
    init_data[1058] = {1'b1,  8'h01};
    init_data[1059] = {1'b1,  8'h03};
    init_data[1060] = {2'b01, 7'h77};
    init_data[1061] = {1'b1,  8'h06};
    init_data[1062] = {1'b1,  8'h14};
    init_data[1063] = {2'b01, 7'h77};
    init_data[1064] = {1'b1,  8'h01};
    init_data[1065] = {1'b1,  8'h03};
    init_data[1066] = {2'b01, 7'h77};
    init_data[1067] = {1'b1,  8'h07};
    init_data[1068] = {1'b1,  8'h00};
    init_data[1069] = {2'b01, 7'h77};
    init_data[1070] = {1'b1,  8'h01};
    init_data[1071] = {1'b1,  8'h03};
    init_data[1072] = {2'b01, 7'h77};
    init_data[1073] = {1'b1,  8'h08};
    init_data[1074] = {1'b1,  8'h00};
    init_data[1075] = {2'b01, 7'h77};
    init_data[1076] = {1'b1,  8'h01};
    init_data[1077] = {1'b1,  8'h03};
    init_data[1078] = {2'b01, 7'h77};
    init_data[1079] = {1'b1,  8'h09};
    init_data[1080] = {1'b1,  8'h00};
    init_data[1081] = {2'b01, 7'h77};
    init_data[1082] = {1'b1,  8'h01};
    init_data[1083] = {1'b1,  8'h03};
    init_data[1084] = {2'b01, 7'h77};
    init_data[1085] = {1'b1,  8'h0A};
    init_data[1086] = {1'b1,  8'h00};
    init_data[1087] = {2'b01, 7'h77};
    init_data[1088] = {1'b1,  8'h01};
    init_data[1089] = {1'b1,  8'h03};
    init_data[1090] = {2'b01, 7'h77};
    init_data[1091] = {1'b1,  8'h0B};
    init_data[1092] = {1'b1,  8'h80};
    init_data[1093] = {2'b01, 7'h77};
    init_data[1094] = {1'b1,  8'h01};
    init_data[1095] = {1'b1,  8'h03};
    init_data[1096] = {2'b01, 7'h77};
    init_data[1097] = {1'b1,  8'h0C};
    init_data[1098] = {1'b1,  8'h00};
    init_data[1099] = {2'b01, 7'h77};
    init_data[1100] = {1'b1,  8'h01};
    init_data[1101] = {1'b1,  8'h03};
    init_data[1102] = {2'b01, 7'h77};
    init_data[1103] = {1'b1,  8'h0D};
    init_data[1104] = {1'b1,  8'h00};
    init_data[1105] = {2'b01, 7'h77};
    init_data[1106] = {1'b1,  8'h01};
    init_data[1107] = {1'b1,  8'h03};
    init_data[1108] = {2'b01, 7'h77};
    init_data[1109] = {1'b1,  8'h0E};
    init_data[1110] = {1'b1,  8'h00};
    init_data[1111] = {2'b01, 7'h77};
    init_data[1112] = {1'b1,  8'h01};
    init_data[1113] = {1'b1,  8'h03};
    init_data[1114] = {2'b01, 7'h77};
    init_data[1115] = {1'b1,  8'h0F};
    init_data[1116] = {1'b1,  8'h00};
    init_data[1117] = {2'b01, 7'h77};
    init_data[1118] = {1'b1,  8'h01};
    init_data[1119] = {1'b1,  8'h03};
    init_data[1120] = {2'b01, 7'h77};
    init_data[1121] = {1'b1,  8'h10};
    init_data[1122] = {1'b1,  8'h00};
    init_data[1123] = {2'b01, 7'h77};
    init_data[1124] = {1'b1,  8'h01};
    init_data[1125] = {1'b1,  8'h03};
    init_data[1126] = {2'b01, 7'h77};
    init_data[1127] = {1'b1,  8'h11};
    init_data[1128] = {1'b1,  8'h00};
    init_data[1129] = {2'b01, 7'h77};
    init_data[1130] = {1'b1,  8'h01};
    init_data[1131] = {1'b1,  8'h03};
    init_data[1132] = {2'b01, 7'h77};
    init_data[1133] = {1'b1,  8'h12};
    init_data[1134] = {1'b1,  8'h00};
    init_data[1135] = {2'b01, 7'h77};
    init_data[1136] = {1'b1,  8'h01};
    init_data[1137] = {1'b1,  8'h03};
    init_data[1138] = {2'b01, 7'h77};
    init_data[1139] = {1'b1,  8'h13};
    init_data[1140] = {1'b1,  8'h00};
    init_data[1141] = {2'b01, 7'h77};
    init_data[1142] = {1'b1,  8'h01};
    init_data[1143] = {1'b1,  8'h03};
    init_data[1144] = {2'b01, 7'h77};
    init_data[1145] = {1'b1,  8'h14};
    init_data[1146] = {1'b1,  8'h00};
    init_data[1147] = {2'b01, 7'h77};
    init_data[1148] = {1'b1,  8'h01};
    init_data[1149] = {1'b1,  8'h03};
    init_data[1150] = {2'b01, 7'h77};
    init_data[1151] = {1'b1,  8'h15};
    init_data[1152] = {1'b1,  8'h00};
    init_data[1153] = {2'b01, 7'h77};
    init_data[1154] = {1'b1,  8'h01};
    init_data[1155] = {1'b1,  8'h03};
    init_data[1156] = {2'b01, 7'h77};
    init_data[1157] = {1'b1,  8'h16};
    init_data[1158] = {1'b1,  8'h00};
    init_data[1159] = {2'b01, 7'h77};
    init_data[1160] = {1'b1,  8'h01};
    init_data[1161] = {1'b1,  8'h03};
    init_data[1162] = {2'b01, 7'h77};
    init_data[1163] = {1'b1,  8'h17};
    init_data[1164] = {1'b1,  8'h00};
    init_data[1165] = {2'b01, 7'h77};
    init_data[1166] = {1'b1,  8'h01};
    init_data[1167] = {1'b1,  8'h03};
    init_data[1168] = {2'b01, 7'h77};
    init_data[1169] = {1'b1,  8'h18};
    init_data[1170] = {1'b1,  8'h00};
    init_data[1171] = {2'b01, 7'h77};
    init_data[1172] = {1'b1,  8'h01};
    init_data[1173] = {1'b1,  8'h03};
    init_data[1174] = {2'b01, 7'h77};
    init_data[1175] = {1'b1,  8'h19};
    init_data[1176] = {1'b1,  8'h00};
    init_data[1177] = {2'b01, 7'h77};
    init_data[1178] = {1'b1,  8'h01};
    init_data[1179] = {1'b1,  8'h03};
    init_data[1180] = {2'b01, 7'h77};
    init_data[1181] = {1'b1,  8'h1A};
    init_data[1182] = {1'b1,  8'h00};
    init_data[1183] = {2'b01, 7'h77};
    init_data[1184] = {1'b1,  8'h01};
    init_data[1185] = {1'b1,  8'h03};
    init_data[1186] = {2'b01, 7'h77};
    init_data[1187] = {1'b1,  8'h1B};
    init_data[1188] = {1'b1,  8'h00};
    init_data[1189] = {2'b01, 7'h77};
    init_data[1190] = {1'b1,  8'h01};
    init_data[1191] = {1'b1,  8'h03};
    init_data[1192] = {2'b01, 7'h77};
    init_data[1193] = {1'b1,  8'h1C};
    init_data[1194] = {1'b1,  8'h00};
    init_data[1195] = {2'b01, 7'h77};
    init_data[1196] = {1'b1,  8'h01};
    init_data[1197] = {1'b1,  8'h03};
    init_data[1198] = {2'b01, 7'h77};
    init_data[1199] = {1'b1,  8'h1D};
    init_data[1200] = {1'b1,  8'h00};
    init_data[1201] = {2'b01, 7'h77};
    init_data[1202] = {1'b1,  8'h01};
    init_data[1203] = {1'b1,  8'h03};
    init_data[1204] = {2'b01, 7'h77};
    init_data[1205] = {1'b1,  8'h1E};
    init_data[1206] = {1'b1,  8'h00};
    init_data[1207] = {2'b01, 7'h77};
    init_data[1208] = {1'b1,  8'h01};
    init_data[1209] = {1'b1,  8'h03};
    init_data[1210] = {2'b01, 7'h77};
    init_data[1211] = {1'b1,  8'h1F};
    init_data[1212] = {1'b1,  8'h00};
    init_data[1213] = {2'b01, 7'h77};
    init_data[1214] = {1'b1,  8'h01};
    init_data[1215] = {1'b1,  8'h03};
    init_data[1216] = {2'b01, 7'h77};
    init_data[1217] = {1'b1,  8'h20};
    init_data[1218] = {1'b1,  8'h00};
    init_data[1219] = {2'b01, 7'h77};
    init_data[1220] = {1'b1,  8'h01};
    init_data[1221] = {1'b1,  8'h03};
    init_data[1222] = {2'b01, 7'h77};
    init_data[1223] = {1'b1,  8'h21};
    init_data[1224] = {1'b1,  8'h00};
    init_data[1225] = {2'b01, 7'h77};
    init_data[1226] = {1'b1,  8'h01};
    init_data[1227] = {1'b1,  8'h03};
    init_data[1228] = {2'b01, 7'h77};
    init_data[1229] = {1'b1,  8'h22};
    init_data[1230] = {1'b1,  8'h00};
    init_data[1231] = {2'b01, 7'h77};
    init_data[1232] = {1'b1,  8'h01};
    init_data[1233] = {1'b1,  8'h03};
    init_data[1234] = {2'b01, 7'h77};
    init_data[1235] = {1'b1,  8'h23};
    init_data[1236] = {1'b1,  8'h00};
    init_data[1237] = {2'b01, 7'h77};
    init_data[1238] = {1'b1,  8'h01};
    init_data[1239] = {1'b1,  8'h03};
    init_data[1240] = {2'b01, 7'h77};
    init_data[1241] = {1'b1,  8'h24};
    init_data[1242] = {1'b1,  8'h00};
    init_data[1243] = {2'b01, 7'h77};
    init_data[1244] = {1'b1,  8'h01};
    init_data[1245] = {1'b1,  8'h03};
    init_data[1246] = {2'b01, 7'h77};
    init_data[1247] = {1'b1,  8'h25};
    init_data[1248] = {1'b1,  8'h00};
    init_data[1249] = {2'b01, 7'h77};
    init_data[1250] = {1'b1,  8'h01};
    init_data[1251] = {1'b1,  8'h03};
    init_data[1252] = {2'b01, 7'h77};
    init_data[1253] = {1'b1,  8'h26};
    init_data[1254] = {1'b1,  8'h00};
    init_data[1255] = {2'b01, 7'h77};
    init_data[1256] = {1'b1,  8'h01};
    init_data[1257] = {1'b1,  8'h03};
    init_data[1258] = {2'b01, 7'h77};
    init_data[1259] = {1'b1,  8'h27};
    init_data[1260] = {1'b1,  8'h00};
    init_data[1261] = {2'b01, 7'h77};
    init_data[1262] = {1'b1,  8'h01};
    init_data[1263] = {1'b1,  8'h03};
    init_data[1264] = {2'b01, 7'h77};
    init_data[1265] = {1'b1,  8'h28};
    init_data[1266] = {1'b1,  8'h00};
    init_data[1267] = {2'b01, 7'h77};
    init_data[1268] = {1'b1,  8'h01};
    init_data[1269] = {1'b1,  8'h03};
    init_data[1270] = {2'b01, 7'h77};
    init_data[1271] = {1'b1,  8'h29};
    init_data[1272] = {1'b1,  8'h00};
    init_data[1273] = {2'b01, 7'h77};
    init_data[1274] = {1'b1,  8'h01};
    init_data[1275] = {1'b1,  8'h03};
    init_data[1276] = {2'b01, 7'h77};
    init_data[1277] = {1'b1,  8'h2A};
    init_data[1278] = {1'b1,  8'h00};
    init_data[1279] = {2'b01, 7'h77};
    init_data[1280] = {1'b1,  8'h01};
    init_data[1281] = {1'b1,  8'h03};
    init_data[1282] = {2'b01, 7'h77};
    init_data[1283] = {1'b1,  8'h2B};
    init_data[1284] = {1'b1,  8'h00};
    init_data[1285] = {2'b01, 7'h77};
    init_data[1286] = {1'b1,  8'h01};
    init_data[1287] = {1'b1,  8'h03};
    init_data[1288] = {2'b01, 7'h77};
    init_data[1289] = {1'b1,  8'h2C};
    init_data[1290] = {1'b1,  8'h00};
    init_data[1291] = {2'b01, 7'h77};
    init_data[1292] = {1'b1,  8'h01};
    init_data[1293] = {1'b1,  8'h03};
    init_data[1294] = {2'b01, 7'h77};
    init_data[1295] = {1'b1,  8'h2D};
    init_data[1296] = {1'b1,  8'h00};
    init_data[1297] = {2'b01, 7'h77};
    init_data[1298] = {1'b1,  8'h01};
    init_data[1299] = {1'b1,  8'h03};
    init_data[1300] = {2'b01, 7'h77};
    init_data[1301] = {1'b1,  8'h2E};
    init_data[1302] = {1'b1,  8'h00};
    init_data[1303] = {2'b01, 7'h77};
    init_data[1304] = {1'b1,  8'h01};
    init_data[1305] = {1'b1,  8'h03};
    init_data[1306] = {2'b01, 7'h77};
    init_data[1307] = {1'b1,  8'h2F};
    init_data[1308] = {1'b1,  8'h00};
    init_data[1309] = {2'b01, 7'h77};
    init_data[1310] = {1'b1,  8'h01};
    init_data[1311] = {1'b1,  8'h03};
    init_data[1312] = {2'b01, 7'h77};
    init_data[1313] = {1'b1,  8'h30};
    init_data[1314] = {1'b1,  8'h00};
    init_data[1315] = {2'b01, 7'h77};
    init_data[1316] = {1'b1,  8'h01};
    init_data[1317] = {1'b1,  8'h03};
    init_data[1318] = {2'b01, 7'h77};
    init_data[1319] = {1'b1,  8'h31};
    init_data[1320] = {1'b1,  8'h00};
    init_data[1321] = {2'b01, 7'h77};
    init_data[1322] = {1'b1,  8'h01};
    init_data[1323] = {1'b1,  8'h03};
    init_data[1324] = {2'b01, 7'h77};
    init_data[1325] = {1'b1,  8'h32};
    init_data[1326] = {1'b1,  8'h00};
    init_data[1327] = {2'b01, 7'h77};
    init_data[1328] = {1'b1,  8'h01};
    init_data[1329] = {1'b1,  8'h03};
    init_data[1330] = {2'b01, 7'h77};
    init_data[1331] = {1'b1,  8'h33};
    init_data[1332] = {1'b1,  8'h00};
    init_data[1333] = {2'b01, 7'h77};
    init_data[1334] = {1'b1,  8'h01};
    init_data[1335] = {1'b1,  8'h03};
    init_data[1336] = {2'b01, 7'h77};
    init_data[1337] = {1'b1,  8'h34};
    init_data[1338] = {1'b1,  8'h00};
    init_data[1339] = {2'b01, 7'h77};
    init_data[1340] = {1'b1,  8'h01};
    init_data[1341] = {1'b1,  8'h03};
    init_data[1342] = {2'b01, 7'h77};
    init_data[1343] = {1'b1,  8'h35};
    init_data[1344] = {1'b1,  8'h00};
    init_data[1345] = {2'b01, 7'h77};
    init_data[1346] = {1'b1,  8'h01};
    init_data[1347] = {1'b1,  8'h03};
    init_data[1348] = {2'b01, 7'h77};
    init_data[1349] = {1'b1,  8'h36};
    init_data[1350] = {1'b1,  8'h00};
    init_data[1351] = {2'b01, 7'h77};
    init_data[1352] = {1'b1,  8'h01};
    init_data[1353] = {1'b1,  8'h03};
    init_data[1354] = {2'b01, 7'h77};
    init_data[1355] = {1'b1,  8'h37};
    init_data[1356] = {1'b1,  8'h00};
    init_data[1357] = {2'b01, 7'h77};
    init_data[1358] = {1'b1,  8'h01};
    init_data[1359] = {1'b1,  8'h03};
    init_data[1360] = {2'b01, 7'h77};
    init_data[1361] = {1'b1,  8'h38};
    init_data[1362] = {1'b1,  8'h00};
    init_data[1363] = {2'b01, 7'h77};
    init_data[1364] = {1'b1,  8'h01};
    init_data[1365] = {1'b1,  8'h03};
    init_data[1366] = {2'b01, 7'h77};
    init_data[1367] = {1'b1,  8'h39};
    init_data[1368] = {1'b1,  8'h1F};
    init_data[1369] = {2'b01, 7'h77};
    init_data[1370] = {1'b1,  8'h01};
    init_data[1371] = {1'b1,  8'h03};
    init_data[1372] = {2'b01, 7'h77};
    init_data[1373] = {1'b1,  8'h3B};
    init_data[1374] = {1'b1,  8'h00};
    init_data[1375] = {2'b01, 7'h77};
    init_data[1376] = {1'b1,  8'h01};
    init_data[1377] = {1'b1,  8'h03};
    init_data[1378] = {2'b01, 7'h77};
    init_data[1379] = {1'b1,  8'h3C};
    init_data[1380] = {1'b1,  8'h00};
    init_data[1381] = {2'b01, 7'h77};
    init_data[1382] = {1'b1,  8'h01};
    init_data[1383] = {1'b1,  8'h03};
    init_data[1384] = {2'b01, 7'h77};
    init_data[1385] = {1'b1,  8'h3D};
    init_data[1386] = {1'b1,  8'h00};
    init_data[1387] = {2'b01, 7'h77};
    init_data[1388] = {1'b1,  8'h01};
    init_data[1389] = {1'b1,  8'h03};
    init_data[1390] = {2'b01, 7'h77};
    init_data[1391] = {1'b1,  8'h3E};
    init_data[1392] = {1'b1,  8'h00};
    init_data[1393] = {2'b01, 7'h77};
    init_data[1394] = {1'b1,  8'h01};
    init_data[1395] = {1'b1,  8'h03};
    init_data[1396] = {2'b01, 7'h77};
    init_data[1397] = {1'b1,  8'h3F};
    init_data[1398] = {1'b1,  8'h00};
    init_data[1399] = {2'b01, 7'h77};
    init_data[1400] = {1'b1,  8'h01};
    init_data[1401] = {1'b1,  8'h03};
    init_data[1402] = {2'b01, 7'h77};
    init_data[1403] = {1'b1,  8'h40};
    init_data[1404] = {1'b1,  8'h00};
    init_data[1405] = {2'b01, 7'h77};
    init_data[1406] = {1'b1,  8'h01};
    init_data[1407] = {1'b1,  8'h03};
    init_data[1408] = {2'b01, 7'h77};
    init_data[1409] = {1'b1,  8'h41};
    init_data[1410] = {1'b1,  8'h00};
    init_data[1411] = {2'b01, 7'h77};
    init_data[1412] = {1'b1,  8'h01};
    init_data[1413] = {1'b1,  8'h03};
    init_data[1414] = {2'b01, 7'h77};
    init_data[1415] = {1'b1,  8'h42};
    init_data[1416] = {1'b1,  8'h00};
    init_data[1417] = {2'b01, 7'h77};
    init_data[1418] = {1'b1,  8'h01};
    init_data[1419] = {1'b1,  8'h03};
    init_data[1420] = {2'b01, 7'h77};
    init_data[1421] = {1'b1,  8'h43};
    init_data[1422] = {1'b1,  8'h00};
    init_data[1423] = {2'b01, 7'h77};
    init_data[1424] = {1'b1,  8'h01};
    init_data[1425] = {1'b1,  8'h03};
    init_data[1426] = {2'b01, 7'h77};
    init_data[1427] = {1'b1,  8'h44};
    init_data[1428] = {1'b1,  8'h00};
    init_data[1429] = {2'b01, 7'h77};
    init_data[1430] = {1'b1,  8'h01};
    init_data[1431] = {1'b1,  8'h03};
    init_data[1432] = {2'b01, 7'h77};
    init_data[1433] = {1'b1,  8'h45};
    init_data[1434] = {1'b1,  8'h00};
    init_data[1435] = {2'b01, 7'h77};
    init_data[1436] = {1'b1,  8'h01};
    init_data[1437] = {1'b1,  8'h03};
    init_data[1438] = {2'b01, 7'h77};
    init_data[1439] = {1'b1,  8'h46};
    init_data[1440] = {1'b1,  8'h00};
    init_data[1441] = {2'b01, 7'h77};
    init_data[1442] = {1'b1,  8'h01};
    init_data[1443] = {1'b1,  8'h03};
    init_data[1444] = {2'b01, 7'h77};
    init_data[1445] = {1'b1,  8'h47};
    init_data[1446] = {1'b1,  8'h00};
    init_data[1447] = {2'b01, 7'h77};
    init_data[1448] = {1'b1,  8'h01};
    init_data[1449] = {1'b1,  8'h03};
    init_data[1450] = {2'b01, 7'h77};
    init_data[1451] = {1'b1,  8'h48};
    init_data[1452] = {1'b1,  8'h00};
    init_data[1453] = {2'b01, 7'h77};
    init_data[1454] = {1'b1,  8'h01};
    init_data[1455] = {1'b1,  8'h03};
    init_data[1456] = {2'b01, 7'h77};
    init_data[1457] = {1'b1,  8'h49};
    init_data[1458] = {1'b1,  8'h00};
    init_data[1459] = {2'b01, 7'h77};
    init_data[1460] = {1'b1,  8'h01};
    init_data[1461] = {1'b1,  8'h03};
    init_data[1462] = {2'b01, 7'h77};
    init_data[1463] = {1'b1,  8'h4A};
    init_data[1464] = {1'b1,  8'h00};
    init_data[1465] = {2'b01, 7'h77};
    init_data[1466] = {1'b1,  8'h01};
    init_data[1467] = {1'b1,  8'h03};
    init_data[1468] = {2'b01, 7'h77};
    init_data[1469] = {1'b1,  8'h4B};
    init_data[1470] = {1'b1,  8'h00};
    init_data[1471] = {2'b01, 7'h77};
    init_data[1472] = {1'b1,  8'h01};
    init_data[1473] = {1'b1,  8'h03};
    init_data[1474] = {2'b01, 7'h77};
    init_data[1475] = {1'b1,  8'h4C};
    init_data[1476] = {1'b1,  8'h00};
    init_data[1477] = {2'b01, 7'h77};
    init_data[1478] = {1'b1,  8'h01};
    init_data[1479] = {1'b1,  8'h03};
    init_data[1480] = {2'b01, 7'h77};
    init_data[1481] = {1'b1,  8'h4D};
    init_data[1482] = {1'b1,  8'h00};
    init_data[1483] = {2'b01, 7'h77};
    init_data[1484] = {1'b1,  8'h01};
    init_data[1485] = {1'b1,  8'h03};
    init_data[1486] = {2'b01, 7'h77};
    init_data[1487] = {1'b1,  8'h4E};
    init_data[1488] = {1'b1,  8'h00};
    init_data[1489] = {2'b01, 7'h77};
    init_data[1490] = {1'b1,  8'h01};
    init_data[1491] = {1'b1,  8'h03};
    init_data[1492] = {2'b01, 7'h77};
    init_data[1493] = {1'b1,  8'h4F};
    init_data[1494] = {1'b1,  8'h00};
    init_data[1495] = {2'b01, 7'h77};
    init_data[1496] = {1'b1,  8'h01};
    init_data[1497] = {1'b1,  8'h03};
    init_data[1498] = {2'b01, 7'h77};
    init_data[1499] = {1'b1,  8'h50};
    init_data[1500] = {1'b1,  8'h00};
    init_data[1501] = {2'b01, 7'h77};
    init_data[1502] = {1'b1,  8'h01};
    init_data[1503] = {1'b1,  8'h03};
    init_data[1504] = {2'b01, 7'h77};
    init_data[1505] = {1'b1,  8'h51};
    init_data[1506] = {1'b1,  8'h00};
    init_data[1507] = {2'b01, 7'h77};
    init_data[1508] = {1'b1,  8'h01};
    init_data[1509] = {1'b1,  8'h03};
    init_data[1510] = {2'b01, 7'h77};
    init_data[1511] = {1'b1,  8'h52};
    init_data[1512] = {1'b1,  8'h00};
    init_data[1513] = {2'b01, 7'h77};
    init_data[1514] = {1'b1,  8'h01};
    init_data[1515] = {1'b1,  8'h03};
    init_data[1516] = {2'b01, 7'h77};
    init_data[1517] = {1'b1,  8'h53};
    init_data[1518] = {1'b1,  8'h00};
    init_data[1519] = {2'b01, 7'h77};
    init_data[1520] = {1'b1,  8'h01};
    init_data[1521] = {1'b1,  8'h03};
    init_data[1522] = {2'b01, 7'h77};
    init_data[1523] = {1'b1,  8'h54};
    init_data[1524] = {1'b1,  8'h00};
    init_data[1525] = {2'b01, 7'h77};
    init_data[1526] = {1'b1,  8'h01};
    init_data[1527] = {1'b1,  8'h03};
    init_data[1528] = {2'b01, 7'h77};
    init_data[1529] = {1'b1,  8'h55};
    init_data[1530] = {1'b1,  8'h00};
    init_data[1531] = {2'b01, 7'h77};
    init_data[1532] = {1'b1,  8'h01};
    init_data[1533] = {1'b1,  8'h03};
    init_data[1534] = {2'b01, 7'h77};
    init_data[1535] = {1'b1,  8'h56};
    init_data[1536] = {1'b1,  8'h00};
    init_data[1537] = {2'b01, 7'h77};
    init_data[1538] = {1'b1,  8'h01};
    init_data[1539] = {1'b1,  8'h03};
    init_data[1540] = {2'b01, 7'h77};
    init_data[1541] = {1'b1,  8'h57};
    init_data[1542] = {1'b1,  8'h00};
    init_data[1543] = {2'b01, 7'h77};
    init_data[1544] = {1'b1,  8'h01};
    init_data[1545] = {1'b1,  8'h03};
    init_data[1546] = {2'b01, 7'h77};
    init_data[1547] = {1'b1,  8'h58};
    init_data[1548] = {1'b1,  8'h00};
    init_data[1549] = {2'b01, 7'h77};
    init_data[1550] = {1'b1,  8'h01};
    init_data[1551] = {1'b1,  8'h03};
    init_data[1552] = {2'b01, 7'h77};
    init_data[1553] = {1'b1,  8'h59};
    init_data[1554] = {1'b1,  8'h00};
    init_data[1555] = {2'b01, 7'h77};
    init_data[1556] = {1'b1,  8'h01};
    init_data[1557] = {1'b1,  8'h03};
    init_data[1558] = {2'b01, 7'h77};
    init_data[1559] = {1'b1,  8'h5A};
    init_data[1560] = {1'b1,  8'h00};
    init_data[1561] = {2'b01, 7'h77};
    init_data[1562] = {1'b1,  8'h01};
    init_data[1563] = {1'b1,  8'h03};
    init_data[1564] = {2'b01, 7'h77};
    init_data[1565] = {1'b1,  8'h5B};
    init_data[1566] = {1'b1,  8'h00};
    init_data[1567] = {2'b01, 7'h77};
    init_data[1568] = {1'b1,  8'h01};
    init_data[1569] = {1'b1,  8'h03};
    init_data[1570] = {2'b01, 7'h77};
    init_data[1571] = {1'b1,  8'h5C};
    init_data[1572] = {1'b1,  8'h00};
    init_data[1573] = {2'b01, 7'h77};
    init_data[1574] = {1'b1,  8'h01};
    init_data[1575] = {1'b1,  8'h03};
    init_data[1576] = {2'b01, 7'h77};
    init_data[1577] = {1'b1,  8'h5D};
    init_data[1578] = {1'b1,  8'h00};
    init_data[1579] = {2'b01, 7'h77};
    init_data[1580] = {1'b1,  8'h01};
    init_data[1581] = {1'b1,  8'h03};
    init_data[1582] = {2'b01, 7'h77};
    init_data[1583] = {1'b1,  8'h5E};
    init_data[1584] = {1'b1,  8'h00};
    init_data[1585] = {2'b01, 7'h77};
    init_data[1586] = {1'b1,  8'h01};
    init_data[1587] = {1'b1,  8'h03};
    init_data[1588] = {2'b01, 7'h77};
    init_data[1589] = {1'b1,  8'h5F};
    init_data[1590] = {1'b1,  8'h00};
    init_data[1591] = {2'b01, 7'h77};
    init_data[1592] = {1'b1,  8'h01};
    init_data[1593] = {1'b1,  8'h03};
    init_data[1594] = {2'b01, 7'h77};
    init_data[1595] = {1'b1,  8'h60};
    init_data[1596] = {1'b1,  8'h00};
    init_data[1597] = {2'b01, 7'h77};
    init_data[1598] = {1'b1,  8'h01};
    init_data[1599] = {1'b1,  8'h03};
    init_data[1600] = {2'b01, 7'h77};
    init_data[1601] = {1'b1,  8'h61};
    init_data[1602] = {1'b1,  8'h00};
    init_data[1603] = {2'b01, 7'h77};
    init_data[1604] = {1'b1,  8'h01};
    init_data[1605] = {1'b1,  8'h03};
    init_data[1606] = {2'b01, 7'h77};
    init_data[1607] = {1'b1,  8'h62};
    init_data[1608] = {1'b1,  8'h00};
    init_data[1609] = {2'b01, 7'h77};
    init_data[1610] = {1'b1,  8'h01};
    init_data[1611] = {1'b1,  8'h08};
    init_data[1612] = {2'b01, 7'h77};
    init_data[1613] = {1'b1,  8'h02};
    init_data[1614] = {1'b1,  8'h00};
    init_data[1615] = {2'b01, 7'h77};
    init_data[1616] = {1'b1,  8'h01};
    init_data[1617] = {1'b1,  8'h08};
    init_data[1618] = {2'b01, 7'h77};
    init_data[1619] = {1'b1,  8'h03};
    init_data[1620] = {1'b1,  8'h00};
    init_data[1621] = {2'b01, 7'h77};
    init_data[1622] = {1'b1,  8'h01};
    init_data[1623] = {1'b1,  8'h08};
    init_data[1624] = {2'b01, 7'h77};
    init_data[1625] = {1'b1,  8'h04};
    init_data[1626] = {1'b1,  8'h00};
    init_data[1627] = {2'b01, 7'h77};
    init_data[1628] = {1'b1,  8'h01};
    init_data[1629] = {1'b1,  8'h08};
    init_data[1630] = {2'b01, 7'h77};
    init_data[1631] = {1'b1,  8'h05};
    init_data[1632] = {1'b1,  8'h00};
    init_data[1633] = {2'b01, 7'h77};
    init_data[1634] = {1'b1,  8'h01};
    init_data[1635] = {1'b1,  8'h08};
    init_data[1636] = {2'b01, 7'h77};
    init_data[1637] = {1'b1,  8'h06};
    init_data[1638] = {1'b1,  8'h00};
    init_data[1639] = {2'b01, 7'h77};
    init_data[1640] = {1'b1,  8'h01};
    init_data[1641] = {1'b1,  8'h08};
    init_data[1642] = {2'b01, 7'h77};
    init_data[1643] = {1'b1,  8'h07};
    init_data[1644] = {1'b1,  8'h00};
    init_data[1645] = {2'b01, 7'h77};
    init_data[1646] = {1'b1,  8'h01};
    init_data[1647] = {1'b1,  8'h08};
    init_data[1648] = {2'b01, 7'h77};
    init_data[1649] = {1'b1,  8'h08};
    init_data[1650] = {1'b1,  8'h00};
    init_data[1651] = {2'b01, 7'h77};
    init_data[1652] = {1'b1,  8'h01};
    init_data[1653] = {1'b1,  8'h08};
    init_data[1654] = {2'b01, 7'h77};
    init_data[1655] = {1'b1,  8'h09};
    init_data[1656] = {1'b1,  8'h00};
    init_data[1657] = {2'b01, 7'h77};
    init_data[1658] = {1'b1,  8'h01};
    init_data[1659] = {1'b1,  8'h08};
    init_data[1660] = {2'b01, 7'h77};
    init_data[1661] = {1'b1,  8'h0A};
    init_data[1662] = {1'b1,  8'h00};
    init_data[1663] = {2'b01, 7'h77};
    init_data[1664] = {1'b1,  8'h01};
    init_data[1665] = {1'b1,  8'h08};
    init_data[1666] = {2'b01, 7'h77};
    init_data[1667] = {1'b1,  8'h0B};
    init_data[1668] = {1'b1,  8'h00};
    init_data[1669] = {2'b01, 7'h77};
    init_data[1670] = {1'b1,  8'h01};
    init_data[1671] = {1'b1,  8'h08};
    init_data[1672] = {2'b01, 7'h77};
    init_data[1673] = {1'b1,  8'h0C};
    init_data[1674] = {1'b1,  8'h00};
    init_data[1675] = {2'b01, 7'h77};
    init_data[1676] = {1'b1,  8'h01};
    init_data[1677] = {1'b1,  8'h08};
    init_data[1678] = {2'b01, 7'h77};
    init_data[1679] = {1'b1,  8'h0D};
    init_data[1680] = {1'b1,  8'h00};
    init_data[1681] = {2'b01, 7'h77};
    init_data[1682] = {1'b1,  8'h01};
    init_data[1683] = {1'b1,  8'h08};
    init_data[1684] = {2'b01, 7'h77};
    init_data[1685] = {1'b1,  8'h0E};
    init_data[1686] = {1'b1,  8'h00};
    init_data[1687] = {2'b01, 7'h77};
    init_data[1688] = {1'b1,  8'h01};
    init_data[1689] = {1'b1,  8'h08};
    init_data[1690] = {2'b01, 7'h77};
    init_data[1691] = {1'b1,  8'h0F};
    init_data[1692] = {1'b1,  8'h00};
    init_data[1693] = {2'b01, 7'h77};
    init_data[1694] = {1'b1,  8'h01};
    init_data[1695] = {1'b1,  8'h08};
    init_data[1696] = {2'b01, 7'h77};
    init_data[1697] = {1'b1,  8'h10};
    init_data[1698] = {1'b1,  8'h00};
    init_data[1699] = {2'b01, 7'h77};
    init_data[1700] = {1'b1,  8'h01};
    init_data[1701] = {1'b1,  8'h08};
    init_data[1702] = {2'b01, 7'h77};
    init_data[1703] = {1'b1,  8'h11};
    init_data[1704] = {1'b1,  8'h00};
    init_data[1705] = {2'b01, 7'h77};
    init_data[1706] = {1'b1,  8'h01};
    init_data[1707] = {1'b1,  8'h08};
    init_data[1708] = {2'b01, 7'h77};
    init_data[1709] = {1'b1,  8'h12};
    init_data[1710] = {1'b1,  8'h00};
    init_data[1711] = {2'b01, 7'h77};
    init_data[1712] = {1'b1,  8'h01};
    init_data[1713] = {1'b1,  8'h08};
    init_data[1714] = {2'b01, 7'h77};
    init_data[1715] = {1'b1,  8'h13};
    init_data[1716] = {1'b1,  8'h00};
    init_data[1717] = {2'b01, 7'h77};
    init_data[1718] = {1'b1,  8'h01};
    init_data[1719] = {1'b1,  8'h08};
    init_data[1720] = {2'b01, 7'h77};
    init_data[1721] = {1'b1,  8'h14};
    init_data[1722] = {1'b1,  8'h00};
    init_data[1723] = {2'b01, 7'h77};
    init_data[1724] = {1'b1,  8'h01};
    init_data[1725] = {1'b1,  8'h08};
    init_data[1726] = {2'b01, 7'h77};
    init_data[1727] = {1'b1,  8'h15};
    init_data[1728] = {1'b1,  8'h00};
    init_data[1729] = {2'b01, 7'h77};
    init_data[1730] = {1'b1,  8'h01};
    init_data[1731] = {1'b1,  8'h08};
    init_data[1732] = {2'b01, 7'h77};
    init_data[1733] = {1'b1,  8'h16};
    init_data[1734] = {1'b1,  8'h00};
    init_data[1735] = {2'b01, 7'h77};
    init_data[1736] = {1'b1,  8'h01};
    init_data[1737] = {1'b1,  8'h08};
    init_data[1738] = {2'b01, 7'h77};
    init_data[1739] = {1'b1,  8'h17};
    init_data[1740] = {1'b1,  8'h00};
    init_data[1741] = {2'b01, 7'h77};
    init_data[1742] = {1'b1,  8'h01};
    init_data[1743] = {1'b1,  8'h08};
    init_data[1744] = {2'b01, 7'h77};
    init_data[1745] = {1'b1,  8'h18};
    init_data[1746] = {1'b1,  8'h00};
    init_data[1747] = {2'b01, 7'h77};
    init_data[1748] = {1'b1,  8'h01};
    init_data[1749] = {1'b1,  8'h08};
    init_data[1750] = {2'b01, 7'h77};
    init_data[1751] = {1'b1,  8'h19};
    init_data[1752] = {1'b1,  8'h00};
    init_data[1753] = {2'b01, 7'h77};
    init_data[1754] = {1'b1,  8'h01};
    init_data[1755] = {1'b1,  8'h08};
    init_data[1756] = {2'b01, 7'h77};
    init_data[1757] = {1'b1,  8'h1A};
    init_data[1758] = {1'b1,  8'h00};
    init_data[1759] = {2'b01, 7'h77};
    init_data[1760] = {1'b1,  8'h01};
    init_data[1761] = {1'b1,  8'h08};
    init_data[1762] = {2'b01, 7'h77};
    init_data[1763] = {1'b1,  8'h1B};
    init_data[1764] = {1'b1,  8'h00};
    init_data[1765] = {2'b01, 7'h77};
    init_data[1766] = {1'b1,  8'h01};
    init_data[1767] = {1'b1,  8'h08};
    init_data[1768] = {2'b01, 7'h77};
    init_data[1769] = {1'b1,  8'h1C};
    init_data[1770] = {1'b1,  8'h00};
    init_data[1771] = {2'b01, 7'h77};
    init_data[1772] = {1'b1,  8'h01};
    init_data[1773] = {1'b1,  8'h08};
    init_data[1774] = {2'b01, 7'h77};
    init_data[1775] = {1'b1,  8'h1D};
    init_data[1776] = {1'b1,  8'h00};
    init_data[1777] = {2'b01, 7'h77};
    init_data[1778] = {1'b1,  8'h01};
    init_data[1779] = {1'b1,  8'h08};
    init_data[1780] = {2'b01, 7'h77};
    init_data[1781] = {1'b1,  8'h1E};
    init_data[1782] = {1'b1,  8'h00};
    init_data[1783] = {2'b01, 7'h77};
    init_data[1784] = {1'b1,  8'h01};
    init_data[1785] = {1'b1,  8'h08};
    init_data[1786] = {2'b01, 7'h77};
    init_data[1787] = {1'b1,  8'h1F};
    init_data[1788] = {1'b1,  8'h00};
    init_data[1789] = {2'b01, 7'h77};
    init_data[1790] = {1'b1,  8'h01};
    init_data[1791] = {1'b1,  8'h08};
    init_data[1792] = {2'b01, 7'h77};
    init_data[1793] = {1'b1,  8'h20};
    init_data[1794] = {1'b1,  8'h00};
    init_data[1795] = {2'b01, 7'h77};
    init_data[1796] = {1'b1,  8'h01};
    init_data[1797] = {1'b1,  8'h08};
    init_data[1798] = {2'b01, 7'h77};
    init_data[1799] = {1'b1,  8'h21};
    init_data[1800] = {1'b1,  8'h00};
    init_data[1801] = {2'b01, 7'h77};
    init_data[1802] = {1'b1,  8'h01};
    init_data[1803] = {1'b1,  8'h08};
    init_data[1804] = {2'b01, 7'h77};
    init_data[1805] = {1'b1,  8'h22};
    init_data[1806] = {1'b1,  8'h00};
    init_data[1807] = {2'b01, 7'h77};
    init_data[1808] = {1'b1,  8'h01};
    init_data[1809] = {1'b1,  8'h08};
    init_data[1810] = {2'b01, 7'h77};
    init_data[1811] = {1'b1,  8'h23};
    init_data[1812] = {1'b1,  8'h00};
    init_data[1813] = {2'b01, 7'h77};
    init_data[1814] = {1'b1,  8'h01};
    init_data[1815] = {1'b1,  8'h08};
    init_data[1816] = {2'b01, 7'h77};
    init_data[1817] = {1'b1,  8'h24};
    init_data[1818] = {1'b1,  8'h00};
    init_data[1819] = {2'b01, 7'h77};
    init_data[1820] = {1'b1,  8'h01};
    init_data[1821] = {1'b1,  8'h08};
    init_data[1822] = {2'b01, 7'h77};
    init_data[1823] = {1'b1,  8'h25};
    init_data[1824] = {1'b1,  8'h00};
    init_data[1825] = {2'b01, 7'h77};
    init_data[1826] = {1'b1,  8'h01};
    init_data[1827] = {1'b1,  8'h08};
    init_data[1828] = {2'b01, 7'h77};
    init_data[1829] = {1'b1,  8'h26};
    init_data[1830] = {1'b1,  8'h00};
    init_data[1831] = {2'b01, 7'h77};
    init_data[1832] = {1'b1,  8'h01};
    init_data[1833] = {1'b1,  8'h08};
    init_data[1834] = {2'b01, 7'h77};
    init_data[1835] = {1'b1,  8'h27};
    init_data[1836] = {1'b1,  8'h00};
    init_data[1837] = {2'b01, 7'h77};
    init_data[1838] = {1'b1,  8'h01};
    init_data[1839] = {1'b1,  8'h08};
    init_data[1840] = {2'b01, 7'h77};
    init_data[1841] = {1'b1,  8'h28};
    init_data[1842] = {1'b1,  8'h00};
    init_data[1843] = {2'b01, 7'h77};
    init_data[1844] = {1'b1,  8'h01};
    init_data[1845] = {1'b1,  8'h08};
    init_data[1846] = {2'b01, 7'h77};
    init_data[1847] = {1'b1,  8'h29};
    init_data[1848] = {1'b1,  8'h00};
    init_data[1849] = {2'b01, 7'h77};
    init_data[1850] = {1'b1,  8'h01};
    init_data[1851] = {1'b1,  8'h08};
    init_data[1852] = {2'b01, 7'h77};
    init_data[1853] = {1'b1,  8'h2A};
    init_data[1854] = {1'b1,  8'h00};
    init_data[1855] = {2'b01, 7'h77};
    init_data[1856] = {1'b1,  8'h01};
    init_data[1857] = {1'b1,  8'h08};
    init_data[1858] = {2'b01, 7'h77};
    init_data[1859] = {1'b1,  8'h2B};
    init_data[1860] = {1'b1,  8'h00};
    init_data[1861] = {2'b01, 7'h77};
    init_data[1862] = {1'b1,  8'h01};
    init_data[1863] = {1'b1,  8'h08};
    init_data[1864] = {2'b01, 7'h77};
    init_data[1865] = {1'b1,  8'h2C};
    init_data[1866] = {1'b1,  8'h00};
    init_data[1867] = {2'b01, 7'h77};
    init_data[1868] = {1'b1,  8'h01};
    init_data[1869] = {1'b1,  8'h08};
    init_data[1870] = {2'b01, 7'h77};
    init_data[1871] = {1'b1,  8'h2D};
    init_data[1872] = {1'b1,  8'h00};
    init_data[1873] = {2'b01, 7'h77};
    init_data[1874] = {1'b1,  8'h01};
    init_data[1875] = {1'b1,  8'h08};
    init_data[1876] = {2'b01, 7'h77};
    init_data[1877] = {1'b1,  8'h2E};
    init_data[1878] = {1'b1,  8'h00};
    init_data[1879] = {2'b01, 7'h77};
    init_data[1880] = {1'b1,  8'h01};
    init_data[1881] = {1'b1,  8'h08};
    init_data[1882] = {2'b01, 7'h77};
    init_data[1883] = {1'b1,  8'h2F};
    init_data[1884] = {1'b1,  8'h00};
    init_data[1885] = {2'b01, 7'h77};
    init_data[1886] = {1'b1,  8'h01};
    init_data[1887] = {1'b1,  8'h08};
    init_data[1888] = {2'b01, 7'h77};
    init_data[1889] = {1'b1,  8'h30};
    init_data[1890] = {1'b1,  8'h00};
    init_data[1891] = {2'b01, 7'h77};
    init_data[1892] = {1'b1,  8'h01};
    init_data[1893] = {1'b1,  8'h08};
    init_data[1894] = {2'b01, 7'h77};
    init_data[1895] = {1'b1,  8'h31};
    init_data[1896] = {1'b1,  8'h00};
    init_data[1897] = {2'b01, 7'h77};
    init_data[1898] = {1'b1,  8'h01};
    init_data[1899] = {1'b1,  8'h08};
    init_data[1900] = {2'b01, 7'h77};
    init_data[1901] = {1'b1,  8'h32};
    init_data[1902] = {1'b1,  8'h00};
    init_data[1903] = {2'b01, 7'h77};
    init_data[1904] = {1'b1,  8'h01};
    init_data[1905] = {1'b1,  8'h08};
    init_data[1906] = {2'b01, 7'h77};
    init_data[1907] = {1'b1,  8'h33};
    init_data[1908] = {1'b1,  8'h00};
    init_data[1909] = {2'b01, 7'h77};
    init_data[1910] = {1'b1,  8'h01};
    init_data[1911] = {1'b1,  8'h08};
    init_data[1912] = {2'b01, 7'h77};
    init_data[1913] = {1'b1,  8'h34};
    init_data[1914] = {1'b1,  8'h00};
    init_data[1915] = {2'b01, 7'h77};
    init_data[1916] = {1'b1,  8'h01};
    init_data[1917] = {1'b1,  8'h08};
    init_data[1918] = {2'b01, 7'h77};
    init_data[1919] = {1'b1,  8'h35};
    init_data[1920] = {1'b1,  8'h00};
    init_data[1921] = {2'b01, 7'h77};
    init_data[1922] = {1'b1,  8'h01};
    init_data[1923] = {1'b1,  8'h08};
    init_data[1924] = {2'b01, 7'h77};
    init_data[1925] = {1'b1,  8'h36};
    init_data[1926] = {1'b1,  8'h00};
    init_data[1927] = {2'b01, 7'h77};
    init_data[1928] = {1'b1,  8'h01};
    init_data[1929] = {1'b1,  8'h08};
    init_data[1930] = {2'b01, 7'h77};
    init_data[1931] = {1'b1,  8'h37};
    init_data[1932] = {1'b1,  8'h00};
    init_data[1933] = {2'b01, 7'h77};
    init_data[1934] = {1'b1,  8'h01};
    init_data[1935] = {1'b1,  8'h08};
    init_data[1936] = {2'b01, 7'h77};
    init_data[1937] = {1'b1,  8'h38};
    init_data[1938] = {1'b1,  8'h00};
    init_data[1939] = {2'b01, 7'h77};
    init_data[1940] = {1'b1,  8'h01};
    init_data[1941] = {1'b1,  8'h08};
    init_data[1942] = {2'b01, 7'h77};
    init_data[1943] = {1'b1,  8'h39};
    init_data[1944] = {1'b1,  8'h00};
    init_data[1945] = {2'b01, 7'h77};
    init_data[1946] = {1'b1,  8'h01};
    init_data[1947] = {1'b1,  8'h08};
    init_data[1948] = {2'b01, 7'h77};
    init_data[1949] = {1'b1,  8'h3A};
    init_data[1950] = {1'b1,  8'h00};
    init_data[1951] = {2'b01, 7'h77};
    init_data[1952] = {1'b1,  8'h01};
    init_data[1953] = {1'b1,  8'h08};
    init_data[1954] = {2'b01, 7'h77};
    init_data[1955] = {1'b1,  8'h3B};
    init_data[1956] = {1'b1,  8'h00};
    init_data[1957] = {2'b01, 7'h77};
    init_data[1958] = {1'b1,  8'h01};
    init_data[1959] = {1'b1,  8'h08};
    init_data[1960] = {2'b01, 7'h77};
    init_data[1961] = {1'b1,  8'h3C};
    init_data[1962] = {1'b1,  8'h00};
    init_data[1963] = {2'b01, 7'h77};
    init_data[1964] = {1'b1,  8'h01};
    init_data[1965] = {1'b1,  8'h08};
    init_data[1966] = {2'b01, 7'h77};
    init_data[1967] = {1'b1,  8'h3D};
    init_data[1968] = {1'b1,  8'h00};
    init_data[1969] = {2'b01, 7'h77};
    init_data[1970] = {1'b1,  8'h01};
    init_data[1971] = {1'b1,  8'h08};
    init_data[1972] = {2'b01, 7'h77};
    init_data[1973] = {1'b1,  8'h3E};
    init_data[1974] = {1'b1,  8'h00};
    init_data[1975] = {2'b01, 7'h77};
    init_data[1976] = {1'b1,  8'h01};
    init_data[1977] = {1'b1,  8'h08};
    init_data[1978] = {2'b01, 7'h77};
    init_data[1979] = {1'b1,  8'h3F};
    init_data[1980] = {1'b1,  8'h00};
    init_data[1981] = {2'b01, 7'h77};
    init_data[1982] = {1'b1,  8'h01};
    init_data[1983] = {1'b1,  8'h08};
    init_data[1984] = {2'b01, 7'h77};
    init_data[1985] = {1'b1,  8'h40};
    init_data[1986] = {1'b1,  8'h00};
    init_data[1987] = {2'b01, 7'h77};
    init_data[1988] = {1'b1,  8'h01};
    init_data[1989] = {1'b1,  8'h08};
    init_data[1990] = {2'b01, 7'h77};
    init_data[1991] = {1'b1,  8'h41};
    init_data[1992] = {1'b1,  8'h00};
    init_data[1993] = {2'b01, 7'h77};
    init_data[1994] = {1'b1,  8'h01};
    init_data[1995] = {1'b1,  8'h08};
    init_data[1996] = {2'b01, 7'h77};
    init_data[1997] = {1'b1,  8'h42};
    init_data[1998] = {1'b1,  8'h00};
    init_data[1999] = {2'b01, 7'h77};
    init_data[2000] = {1'b1,  8'h01};
    init_data[2001] = {1'b1,  8'h08};
    init_data[2002] = {2'b01, 7'h77};
    init_data[2003] = {1'b1,  8'h43};
    init_data[2004] = {1'b1,  8'h00};
    init_data[2005] = {2'b01, 7'h77};
    init_data[2006] = {1'b1,  8'h01};
    init_data[2007] = {1'b1,  8'h08};
    init_data[2008] = {2'b01, 7'h77};
    init_data[2009] = {1'b1,  8'h44};
    init_data[2010] = {1'b1,  8'h00};
    init_data[2011] = {2'b01, 7'h77};
    init_data[2012] = {1'b1,  8'h01};
    init_data[2013] = {1'b1,  8'h08};
    init_data[2014] = {2'b01, 7'h77};
    init_data[2015] = {1'b1,  8'h45};
    init_data[2016] = {1'b1,  8'h00};
    init_data[2017] = {2'b01, 7'h77};
    init_data[2018] = {1'b1,  8'h01};
    init_data[2019] = {1'b1,  8'h08};
    init_data[2020] = {2'b01, 7'h77};
    init_data[2021] = {1'b1,  8'h46};
    init_data[2022] = {1'b1,  8'h00};
    init_data[2023] = {2'b01, 7'h77};
    init_data[2024] = {1'b1,  8'h01};
    init_data[2025] = {1'b1,  8'h08};
    init_data[2026] = {2'b01, 7'h77};
    init_data[2027] = {1'b1,  8'h47};
    init_data[2028] = {1'b1,  8'h00};
    init_data[2029] = {2'b01, 7'h77};
    init_data[2030] = {1'b1,  8'h01};
    init_data[2031] = {1'b1,  8'h08};
    init_data[2032] = {2'b01, 7'h77};
    init_data[2033] = {1'b1,  8'h48};
    init_data[2034] = {1'b1,  8'h00};
    init_data[2035] = {2'b01, 7'h77};
    init_data[2036] = {1'b1,  8'h01};
    init_data[2037] = {1'b1,  8'h08};
    init_data[2038] = {2'b01, 7'h77};
    init_data[2039] = {1'b1,  8'h49};
    init_data[2040] = {1'b1,  8'h00};
    init_data[2041] = {2'b01, 7'h77};
    init_data[2042] = {1'b1,  8'h01};
    init_data[2043] = {1'b1,  8'h08};
    init_data[2044] = {2'b01, 7'h77};
    init_data[2045] = {1'b1,  8'h4A};
    init_data[2046] = {1'b1,  8'h00};
    init_data[2047] = {2'b01, 7'h77};
    init_data[2048] = {1'b1,  8'h01};
    init_data[2049] = {1'b1,  8'h08};
    init_data[2050] = {2'b01, 7'h77};
    init_data[2051] = {1'b1,  8'h4B};
    init_data[2052] = {1'b1,  8'h00};
    init_data[2053] = {2'b01, 7'h77};
    init_data[2054] = {1'b1,  8'h01};
    init_data[2055] = {1'b1,  8'h08};
    init_data[2056] = {2'b01, 7'h77};
    init_data[2057] = {1'b1,  8'h4C};
    init_data[2058] = {1'b1,  8'h00};
    init_data[2059] = {2'b01, 7'h77};
    init_data[2060] = {1'b1,  8'h01};
    init_data[2061] = {1'b1,  8'h08};
    init_data[2062] = {2'b01, 7'h77};
    init_data[2063] = {1'b1,  8'h4D};
    init_data[2064] = {1'b1,  8'h00};
    init_data[2065] = {2'b01, 7'h77};
    init_data[2066] = {1'b1,  8'h01};
    init_data[2067] = {1'b1,  8'h08};
    init_data[2068] = {2'b01, 7'h77};
    init_data[2069] = {1'b1,  8'h4E};
    init_data[2070] = {1'b1,  8'h00};
    init_data[2071] = {2'b01, 7'h77};
    init_data[2072] = {1'b1,  8'h01};
    init_data[2073] = {1'b1,  8'h08};
    init_data[2074] = {2'b01, 7'h77};
    init_data[2075] = {1'b1,  8'h4F};
    init_data[2076] = {1'b1,  8'h00};
    init_data[2077] = {2'b01, 7'h77};
    init_data[2078] = {1'b1,  8'h01};
    init_data[2079] = {1'b1,  8'h08};
    init_data[2080] = {2'b01, 7'h77};
    init_data[2081] = {1'b1,  8'h50};
    init_data[2082] = {1'b1,  8'h00};
    init_data[2083] = {2'b01, 7'h77};
    init_data[2084] = {1'b1,  8'h01};
    init_data[2085] = {1'b1,  8'h08};
    init_data[2086] = {2'b01, 7'h77};
    init_data[2087] = {1'b1,  8'h51};
    init_data[2088] = {1'b1,  8'h00};
    init_data[2089] = {2'b01, 7'h77};
    init_data[2090] = {1'b1,  8'h01};
    init_data[2091] = {1'b1,  8'h08};
    init_data[2092] = {2'b01, 7'h77};
    init_data[2093] = {1'b1,  8'h52};
    init_data[2094] = {1'b1,  8'h00};
    init_data[2095] = {2'b01, 7'h77};
    init_data[2096] = {1'b1,  8'h01};
    init_data[2097] = {1'b1,  8'h08};
    init_data[2098] = {2'b01, 7'h77};
    init_data[2099] = {1'b1,  8'h53};
    init_data[2100] = {1'b1,  8'h00};
    init_data[2101] = {2'b01, 7'h77};
    init_data[2102] = {1'b1,  8'h01};
    init_data[2103] = {1'b1,  8'h08};
    init_data[2104] = {2'b01, 7'h77};
    init_data[2105] = {1'b1,  8'h54};
    init_data[2106] = {1'b1,  8'h00};
    init_data[2107] = {2'b01, 7'h77};
    init_data[2108] = {1'b1,  8'h01};
    init_data[2109] = {1'b1,  8'h08};
    init_data[2110] = {2'b01, 7'h77};
    init_data[2111] = {1'b1,  8'h55};
    init_data[2112] = {1'b1,  8'h00};
    init_data[2113] = {2'b01, 7'h77};
    init_data[2114] = {1'b1,  8'h01};
    init_data[2115] = {1'b1,  8'h08};
    init_data[2116] = {2'b01, 7'h77};
    init_data[2117] = {1'b1,  8'h56};
    init_data[2118] = {1'b1,  8'h00};
    init_data[2119] = {2'b01, 7'h77};
    init_data[2120] = {1'b1,  8'h01};
    init_data[2121] = {1'b1,  8'h08};
    init_data[2122] = {2'b01, 7'h77};
    init_data[2123] = {1'b1,  8'h57};
    init_data[2124] = {1'b1,  8'h00};
    init_data[2125] = {2'b01, 7'h77};
    init_data[2126] = {1'b1,  8'h01};
    init_data[2127] = {1'b1,  8'h08};
    init_data[2128] = {2'b01, 7'h77};
    init_data[2129] = {1'b1,  8'h58};
    init_data[2130] = {1'b1,  8'h00};
    init_data[2131] = {2'b01, 7'h77};
    init_data[2132] = {1'b1,  8'h01};
    init_data[2133] = {1'b1,  8'h08};
    init_data[2134] = {2'b01, 7'h77};
    init_data[2135] = {1'b1,  8'h59};
    init_data[2136] = {1'b1,  8'h00};
    init_data[2137] = {2'b01, 7'h77};
    init_data[2138] = {1'b1,  8'h01};
    init_data[2139] = {1'b1,  8'h08};
    init_data[2140] = {2'b01, 7'h77};
    init_data[2141] = {1'b1,  8'h5A};
    init_data[2142] = {1'b1,  8'h00};
    init_data[2143] = {2'b01, 7'h77};
    init_data[2144] = {1'b1,  8'h01};
    init_data[2145] = {1'b1,  8'h08};
    init_data[2146] = {2'b01, 7'h77};
    init_data[2147] = {1'b1,  8'h5B};
    init_data[2148] = {1'b1,  8'h00};
    init_data[2149] = {2'b01, 7'h77};
    init_data[2150] = {1'b1,  8'h01};
    init_data[2151] = {1'b1,  8'h08};
    init_data[2152] = {2'b01, 7'h77};
    init_data[2153] = {1'b1,  8'h5C};
    init_data[2154] = {1'b1,  8'h00};
    init_data[2155] = {2'b01, 7'h77};
    init_data[2156] = {1'b1,  8'h01};
    init_data[2157] = {1'b1,  8'h08};
    init_data[2158] = {2'b01, 7'h77};
    init_data[2159] = {1'b1,  8'h5D};
    init_data[2160] = {1'b1,  8'h00};
    init_data[2161] = {2'b01, 7'h77};
    init_data[2162] = {1'b1,  8'h01};
    init_data[2163] = {1'b1,  8'h08};
    init_data[2164] = {2'b01, 7'h77};
    init_data[2165] = {1'b1,  8'h5E};
    init_data[2166] = {1'b1,  8'h00};
    init_data[2167] = {2'b01, 7'h77};
    init_data[2168] = {1'b1,  8'h01};
    init_data[2169] = {1'b1,  8'h08};
    init_data[2170] = {2'b01, 7'h77};
    init_data[2171] = {1'b1,  8'h5F};
    init_data[2172] = {1'b1,  8'h00};
    init_data[2173] = {2'b01, 7'h77};
    init_data[2174] = {1'b1,  8'h01};
    init_data[2175] = {1'b1,  8'h08};
    init_data[2176] = {2'b01, 7'h77};
    init_data[2177] = {1'b1,  8'h60};
    init_data[2178] = {1'b1,  8'h00};
    init_data[2179] = {2'b01, 7'h77};
    init_data[2180] = {1'b1,  8'h01};
    init_data[2181] = {1'b1,  8'h08};
    init_data[2182] = {2'b01, 7'h77};
    init_data[2183] = {1'b1,  8'h61};
    init_data[2184] = {1'b1,  8'h00};
    init_data[2185] = {2'b01, 7'h77};
    init_data[2186] = {1'b1,  8'h01};
    init_data[2187] = {1'b1,  8'h09};
    init_data[2188] = {2'b01, 7'h77};
    init_data[2189] = {1'b1,  8'h0E};
    init_data[2190] = {1'b1,  8'h00};
    init_data[2191] = {2'b01, 7'h77};
    init_data[2192] = {1'b1,  8'h01};
    init_data[2193] = {1'b1,  8'h09};
    init_data[2194] = {2'b01, 7'h77};
    init_data[2195] = {1'b1,  8'h1C};
    init_data[2196] = {1'b1,  8'h04};
    init_data[2197] = {2'b01, 7'h77};
    init_data[2198] = {1'b1,  8'h01};
    init_data[2199] = {1'b1,  8'h09};
    init_data[2200] = {2'b01, 7'h77};
    init_data[2201] = {1'b1,  8'h43};
    init_data[2202] = {1'b1,  8'h00};
    init_data[2203] = {2'b01, 7'h77};
    init_data[2204] = {1'b1,  8'h01};
    init_data[2205] = {1'b1,  8'h09};
    init_data[2206] = {2'b01, 7'h77};
    init_data[2207] = {1'b1,  8'h49};
    init_data[2208] = {1'b1,  8'h01};
    init_data[2209] = {2'b01, 7'h77};
    init_data[2210] = {1'b1,  8'h01};
    init_data[2211] = {1'b1,  8'h09};
    init_data[2212] = {2'b01, 7'h77};
    init_data[2213] = {1'b1,  8'h4A};
    init_data[2214] = {1'b1,  8'h10};
    init_data[2215] = {2'b01, 7'h77};
    init_data[2216] = {1'b1,  8'h01};
    init_data[2217] = {1'b1,  8'h09};
    init_data[2218] = {2'b01, 7'h77};
    init_data[2219] = {1'b1,  8'h4E};
    init_data[2220] = {1'b1,  8'h49};
    init_data[2221] = {2'b01, 7'h77};
    init_data[2222] = {1'b1,  8'h01};
    init_data[2223] = {1'b1,  8'h09};
    init_data[2224] = {2'b01, 7'h77};
    init_data[2225] = {1'b1,  8'h4F};
    init_data[2226] = {1'b1,  8'h02};
    init_data[2227] = {2'b01, 7'h77};
    init_data[2228] = {1'b1,  8'h01};
    init_data[2229] = {1'b1,  8'h09};
    init_data[2230] = {2'b01, 7'h77};
    init_data[2231] = {1'b1,  8'h5E};
    init_data[2232] = {1'b1,  8'h00};
    init_data[2233] = {2'b01, 7'h77};
    init_data[2234] = {1'b1,  8'h01};
    init_data[2235] = {1'b1,  8'h0A};
    init_data[2236] = {2'b01, 7'h77};
    init_data[2237] = {1'b1,  8'h02};
    init_data[2238] = {1'b1,  8'h00};
    init_data[2239] = {2'b01, 7'h77};
    init_data[2240] = {1'b1,  8'h01};
    init_data[2241] = {1'b1,  8'h0A};
    init_data[2242] = {2'b01, 7'h77};
    init_data[2243] = {1'b1,  8'h03};
    init_data[2244] = {1'b1,  8'h01};
    init_data[2245] = {2'b01, 7'h77};
    init_data[2246] = {1'b1,  8'h01};
    init_data[2247] = {1'b1,  8'h0A};
    init_data[2248] = {2'b01, 7'h77};
    init_data[2249] = {1'b1,  8'h04};
    init_data[2250] = {1'b1,  8'h01};
    init_data[2251] = {2'b01, 7'h77};
    init_data[2252] = {1'b1,  8'h01};
    init_data[2253] = {1'b1,  8'h0A};
    init_data[2254] = {2'b01, 7'h77};
    init_data[2255] = {1'b1,  8'h05};
    init_data[2256] = {1'b1,  8'h01};
    init_data[2257] = {2'b01, 7'h77};
    init_data[2258] = {1'b1,  8'h01};
    init_data[2259] = {1'b1,  8'h0A};
    init_data[2260] = {2'b01, 7'h77};
    init_data[2261] = {1'b1,  8'h14};
    init_data[2262] = {1'b1,  8'h00};
    init_data[2263] = {2'b01, 7'h77};
    init_data[2264] = {1'b1,  8'h01};
    init_data[2265] = {1'b1,  8'h0A};
    init_data[2266] = {2'b01, 7'h77};
    init_data[2267] = {1'b1,  8'h1A};
    init_data[2268] = {1'b1,  8'h00};
    init_data[2269] = {2'b01, 7'h77};
    init_data[2270] = {1'b1,  8'h01};
    init_data[2271] = {1'b1,  8'h0A};
    init_data[2272] = {2'b01, 7'h77};
    init_data[2273] = {1'b1,  8'h20};
    init_data[2274] = {1'b1,  8'h00};
    init_data[2275] = {2'b01, 7'h77};
    init_data[2276] = {1'b1,  8'h01};
    init_data[2277] = {1'b1,  8'h0A};
    init_data[2278] = {2'b01, 7'h77};
    init_data[2279] = {1'b1,  8'h26};
    init_data[2280] = {1'b1,  8'h00};
    init_data[2281] = {2'b01, 7'h77};
    init_data[2282] = {1'b1,  8'h01};
    init_data[2283] = {1'b1,  8'h0A};
    init_data[2284] = {2'b01, 7'h77};
    init_data[2285] = {1'b1,  8'h2C};
    init_data[2286] = {1'b1,  8'h00};
    init_data[2287] = {2'b01, 7'h77};
    init_data[2288] = {1'b1,  8'h01};
    init_data[2289] = {1'b1,  8'h0B};
    init_data[2290] = {2'b01, 7'h77};
    init_data[2291] = {1'b1,  8'h44};
    init_data[2292] = {1'b1,  8'h0F};
    init_data[2293] = {2'b01, 7'h77};
    init_data[2294] = {1'b1,  8'h01};
    init_data[2295] = {1'b1,  8'h0B};
    init_data[2296] = {2'b01, 7'h77};
    init_data[2297] = {1'b1,  8'h4A};
    init_data[2298] = {1'b1,  8'h1E};
    init_data[2299] = {2'b01, 7'h77};
    init_data[2300] = {1'b1,  8'h01};
    init_data[2301] = {1'b1,  8'h0B};
    init_data[2302] = {2'b01, 7'h77};
    init_data[2303] = {1'b1,  8'h57};
    init_data[2304] = {1'b1,  8'hA5};
    init_data[2305] = {2'b01, 7'h77};
    init_data[2306] = {1'b1,  8'h01};
    init_data[2307] = {1'b1,  8'h0B};
    init_data[2308] = {2'b01, 7'h77};
    init_data[2309] = {1'b1,  8'h58};
    init_data[2310] = {1'b1,  8'h00};
    init_data[2311] = {2'b01, 7'h77};
    init_data[2312] = {1'b1,  8'h01};
    init_data[2313] = {1'b1,  8'h00};
    init_data[2314] = {2'b01, 7'h77};
    init_data[2315] = {1'b1,  8'h1C};
    init_data[2316] = {1'b1,  8'h01};
    init_data[2317] = {2'b01, 7'h77};
    init_data[2318] = {1'b1,  8'h01};
    init_data[2319] = {1'b1,  8'h0B};
    init_data[2320] = {2'b01, 7'h77};
    init_data[2321] = {1'b1,  8'h24};
    init_data[2322] = {1'b1,  8'hC3};
    init_data[2323] = {2'b01, 7'h77};
    init_data[2324] = {1'b1,  8'h01};
    init_data[2325] = {1'b1,  8'h0B};
    init_data[2326] = {2'b01, 7'h77};
    init_data[2327] = {1'b1,  8'h25};
    init_data[2328] = {1'b1,  8'h02};
end

localparam [3:0]
    STATE_IDLE = 3'd0,
    STATE_RUN = 3'd1,
    STATE_TABLE_1 = 3'd2,
    STATE_TABLE_2 = 3'd3,
    STATE_TABLE_3 = 3'd4;

reg [4:0] state_reg = STATE_IDLE, state_next;

parameter AW = $clog2(INIT_DATA_LEN);

reg [8:0] init_data_reg = 9'd0;

reg [31:0] delay_counter = 32'd0;

reg [AW-1:0] address_reg = {AW{1'b0}}, address_next;
reg [AW-1:0] address_ptr_reg = {AW{1'b0}}, address_ptr_next;
reg [AW-1:0] data_ptr_reg = {AW{1'b0}}, data_ptr_next;

reg [6:0] cur_address_reg = 7'd0, cur_address_next;

reg [6:0] cmd_address_reg = 7'd0, cmd_address_next;
reg cmd_start_reg = 1'b0, cmd_start_next;
reg cmd_write_reg = 1'b0, cmd_write_next;
reg cmd_stop_reg = 1'b0, cmd_stop_next;
reg cmd_valid_reg = 1'b0, cmd_valid_next;

reg [7:0] data_out_reg = 8'd0, data_out_next;
reg data_out_valid_reg = 1'b0, data_out_valid_next;

reg start_flag_reg = 1'b0, start_flag_next;

reg busy_reg = 1'b0;

assign cmd_address = cmd_address_reg;
assign cmd_start = cmd_start_reg;
assign cmd_read = 1'b0;
assign cmd_write = cmd_write_reg;
assign cmd_write_multiple = 1'b0;
assign cmd_stop = cmd_stop_reg;
assign cmd_valid = cmd_valid_reg;

assign data_out = data_out_reg;
assign data_out_valid = data_out_valid_reg;
assign data_out_last = 1'b1;

assign busy = busy_reg;

always @* begin
    state_next = STATE_IDLE;

    address_next = address_reg;
    address_ptr_next = address_ptr_reg;
    data_ptr_next = data_ptr_reg;

    cur_address_next = cur_address_reg;

    cmd_address_next = cmd_address_reg;
    cmd_start_next = cmd_start_reg & ~(cmd_valid & cmd_ready);
    cmd_write_next = cmd_write_reg & ~(cmd_valid & cmd_ready);
    cmd_stop_next = cmd_stop_reg & ~(cmd_valid & cmd_ready);
    cmd_valid_next = cmd_valid_reg & ~cmd_ready;

    data_out_next = data_out_reg;
    data_out_valid_next = data_out_valid_reg & ~data_out_ready;

    start_flag_next = start_flag_reg;

    if (cmd_valid | data_out_valid) begin
        // wait for output registers to clear
        state_next = state_reg;
    end else begin
        case (state_reg)
            STATE_IDLE: begin
                // wait for start signal
                if (~start_flag_reg & start) begin
                    address_next = {AW{1'b0}};
                    start_flag_next = 1'b1;
                    state_next = STATE_RUN;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_RUN: begin
                // process commands
                if (init_data_reg[8] == 1'b1) begin
                    // write data
                    cmd_write_next = 1'b1;
                    cmd_stop_next = 1'b0;
                    cmd_valid_next = 1'b1;

                    data_out_next = init_data_reg[7:0];
                    data_out_valid_next = 1'b1;

                    address_next = address_reg + 1;

                    state_next = STATE_RUN;
                end else if (init_data_reg == 9'b111111111) begin
                    //
                    // Delay 300 ms
                    // clk_125mhz
                    // == 37500000 cycles
                    // == 0x23c3460 cycles
                    // 27 bit = 1
                    //
                    if (!delay_counter[27]) begin
                        delay_counter <= delay_counter + 32'd1;
                    end else begin
                        address_next = address_reg + 1;
                    end
                    state_next = STATE_RUN;
                end else if (init_data_reg[8:7] == 2'b01) begin
                    // write address
                    cmd_address_next = init_data_reg[6:0];
                    cmd_start_next = 1'b1;

                    address_next = address_reg + 1;

                    state_next = STATE_RUN;
                end else if (init_data_reg == 9'b001000001) begin
                    // send stop
                    cmd_write_next = 1'b0;
                    cmd_start_next = 1'b0;
                    cmd_stop_next = 1'b1;
                    cmd_valid_next = 1'b1;

                    address_next = address_reg + 1;

                    state_next = STATE_RUN;
                end else if (init_data_reg == 9'b000001001) begin
                    // data table start
                    data_ptr_next = address_reg + 1;
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_1;
                end else if (init_data_reg == 9'd0) begin
                    // stop
                    cmd_start_next = 1'b0;
                    cmd_write_next = 1'b0;
                    cmd_stop_next = 1'b1;
                    cmd_valid_next = 1'b1;

                    state_next = STATE_IDLE;
                end else begin
                    // invalid command, skip
                    address_next = address_reg + 1;
                    state_next = STATE_RUN;
                end
            end
            STATE_TABLE_1: begin
                // find address table start
                if (init_data_reg == 9'b000001000) begin
                    // address table start
                    address_ptr_next = address_reg + 1;
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_2;
                end else if (init_data_reg == 9'b000001001) begin
                    // data table start
                    data_ptr_next = address_reg + 1;
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_1;
                end else if (init_data_reg == 1) begin
                    // exit mode
                    address_next = address_reg + 1;
                    state_next = STATE_RUN;
                end else if (init_data_reg == 9'd0) begin
                    // stop
                    cmd_start_next = 1'b0;
                    cmd_write_next = 1'b0;
                    cmd_stop_next = 1'b1;
                    cmd_valid_next = 1'b1;

                    state_next = STATE_IDLE;
                end else begin
                    // invalid command, skip
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_1;
                end
            end
            STATE_TABLE_2: begin
                // find next address
                if (init_data_reg[8:7] == 2'b01) begin
                    // write address command
                    // store address and move to data table
                    cur_address_next = init_data_reg[6:0];
                    address_ptr_next = address_reg + 1;
                    address_next = data_ptr_reg;
                    state_next = STATE_TABLE_3;
                end else if (init_data_reg == 9'b000001001) begin
                    // data table start
                    data_ptr_next = address_reg + 1;
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_1;
                end else if (init_data_reg == 9'd1) begin
                    // exit mode
                    address_next = address_reg + 1;
                    state_next = STATE_RUN;
                end else if (init_data_reg == 9'd0) begin
                    // stop
                    cmd_start_next = 1'b0;
                    cmd_write_next = 1'b0;
                    cmd_stop_next = 1'b1;
                    cmd_valid_next = 1'b1;

                    state_next = STATE_IDLE;
                end else begin
                    // invalid command, skip
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_2;
                end
            end
            STATE_TABLE_3: begin
                // process data table with selected address
                if (init_data_reg[8] == 1'b1) begin
                    // write data
                    cmd_write_next = 1'b1;
                    cmd_stop_next = 1'b0;
                    cmd_valid_next = 1'b1;

                    data_out_next = init_data_reg[7:0];
                    data_out_valid_next = 1'b1;

                    address_next = address_reg + 1;

                    state_next = STATE_TABLE_3;
                end else if (init_data_reg[8:7] == 2'b01) begin
                    // write address
                    cmd_address_next = init_data_reg[6:0];
                    cmd_start_next = 1'b1;

                    address_next = address_reg + 1;

                    state_next = STATE_TABLE_3;
                end else if (init_data_reg == 9'b000000011) begin
                    // write current address
                    cmd_address_next = cur_address_reg;
                    cmd_start_next = 1'b1;

                    address_next = address_reg + 1;

                    state_next = STATE_TABLE_3;
                end else if (init_data_reg == 9'b001000001) begin
                    // send stop
                    cmd_write_next = 1'b0;
                    cmd_start_next = 1'b0;
                    cmd_stop_next = 1'b1;
                    cmd_valid_next = 1'b1;

                    address_next = address_reg + 1;

                    state_next = STATE_TABLE_3;
                end else if (init_data_reg == 9'b000001001) begin
                    // data table start
                    data_ptr_next = address_reg + 1;
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_1;
                end else if (init_data_reg == 9'b000001000) begin
                    // address table start
                    address_next = address_ptr_reg;
                    state_next = STATE_TABLE_2;
                end else if (init_data_reg == 9'd1) begin
                    // exit mode
                    address_next = address_reg + 1;
                    state_next = STATE_RUN;
                end else if (init_data_reg == 9'd0) begin
                    // stop
                    cmd_start_next = 1'b0;
                    cmd_write_next = 1'b0;
                    cmd_stop_next = 1'b1;
                    cmd_valid_next = 1'b1;

                    state_next = STATE_IDLE;
                end else begin
                    // invalid command, skip
                    address_next = address_reg + 1;
                    state_next = STATE_TABLE_3;
                end
            end
        endcase
    end
end

always @(posedge clk) begin
    if (rst) begin
        state_reg <= STATE_IDLE;

        init_data_reg <= 9'd0;

        address_reg <= {AW{1'b0}};
        address_ptr_reg <= {AW{1'b0}};
        data_ptr_reg <= {AW{1'b0}};

        cur_address_reg <= 7'd0;

        cmd_valid_reg <= 1'b0;

        data_out_valid_reg <= 1'b0;

        start_flag_reg <= 1'b0;

        busy_reg <= 1'b0;
    end else begin
        state_reg <= state_next;

        // read init_data ROM
        init_data_reg <= init_data[address_next];

        address_reg <= address_next;
        address_ptr_reg <= address_ptr_next;
        data_ptr_reg <= data_ptr_next;

        cur_address_reg <= cur_address_next;

        cmd_valid_reg <= cmd_valid_next;

        data_out_valid_reg <= data_out_valid_next;

        start_flag_reg <= start & start_flag_next;

        busy_reg <= (state_reg != STATE_IDLE);
    end

    cmd_address_reg <= cmd_address_next;
    cmd_start_reg <= cmd_start_next;
    cmd_write_reg <= cmd_write_next;
    cmd_stop_reg <= cmd_stop_next;

    data_out_reg <= data_out_next;
end

endmodule
